`include "define.v"

module Image_Classifier ( 
    input clk, 
    input GlobalReset, 
    input Input_Valid,
    input [18:0] Wgt_0_0, // sfix19_En18 
    input [18:0] Wgt_0_1, // sfix19_En18 
    input [18:0] Wgt_0_2, // sfix19_En18 
    input [18:0] Wgt_0_3, // sfix19_En18 
    input [18:0] Wgt_0_4, // sfix19_En18 
    input [18:0] Wgt_0_5, // sfix19_En18 
    input [18:0] Wgt_0_6, // sfix19_En18 
    input [18:0] Wgt_0_7, // sfix19_En18 
    input [18:0] Wgt_0_8, // sfix19_En18 
    input [18:0] Wgt_0_9, // sfix19_En18 
    input [18:0] Wgt_0_10, // sfix19_En18 
    input [18:0] Wgt_0_11, // sfix19_En18 
    input [18:0] Wgt_0_12, // sfix19_En18 
    input [18:0] Wgt_0_13, // sfix19_En18 
    input [18:0] Wgt_0_14, // sfix19_En18 
    input [18:0] Wgt_0_15, // sfix19_En18 
    input [18:0] Wgt_0_16, // sfix19_En18 
    input [18:0] Wgt_0_17, // sfix19_En18 
    input [18:0] Wgt_0_18, // sfix19_En18 
    input [18:0] Wgt_0_19, // sfix19_En18 
    input [18:0] Wgt_0_20, // sfix19_En18 
    input [18:0] Wgt_0_21, // sfix19_En18 
    input [18:0] Wgt_0_22, // sfix19_En18 
    input [18:0] Wgt_0_23, // sfix19_En18 
    input [18:0] Wgt_0_24, // sfix19_En18 
    input [18:0] Wgt_0_25, // sfix19_En18 
    input [18:0] Wgt_0_26, // sfix19_En18 
    input [18:0] Wgt_0_27, // sfix19_En18 
    input [18:0] Wgt_0_28, // sfix19_En18 
    input [18:0] Wgt_0_29, // sfix19_En18 
    input [18:0] Wgt_0_30, // sfix19_En18 
    input [18:0] Wgt_0_31, // sfix19_En18 
    input [18:0] Wgt_0_32, // sfix19_En18 
    input [18:0] Wgt_0_33, // sfix19_En18 
    input [18:0] Wgt_0_34, // sfix19_En18 
    input [18:0] Wgt_0_35, // sfix19_En18 
    input [18:0] Wgt_0_36, // sfix19_En18 
    input [18:0] Wgt_0_37, // sfix19_En18 
    input [18:0] Wgt_0_38, // sfix19_En18 
    input [18:0] Wgt_0_39, // sfix19_En18 
    input [18:0] Wgt_0_40, // sfix19_En18 
    input [18:0] Wgt_0_41, // sfix19_En18 
    input [18:0] Wgt_0_42, // sfix19_En18 
    input [18:0] Wgt_0_43, // sfix19_En18 
    input [18:0] Wgt_0_44, // sfix19_En18 
    input [18:0] Wgt_0_45, // sfix19_En18 
    input [18:0] Wgt_0_46, // sfix19_En18 
    input [18:0] Wgt_0_47, // sfix19_En18 
    input [18:0] Wgt_0_48, // sfix19_En18 
    input [18:0] Wgt_0_49, // sfix19_En18 
    input [18:0] Wgt_0_50, // sfix19_En18 
    input [18:0] Wgt_0_51, // sfix19_En18 
    input [18:0] Wgt_0_52, // sfix19_En18 
    input [18:0] Wgt_0_53, // sfix19_En18 
    input [18:0] Wgt_0_54, // sfix19_En18 
    input [18:0] Wgt_0_55, // sfix19_En18 
    input [18:0] Wgt_0_56, // sfix19_En18 
    input [18:0] Wgt_0_57, // sfix19_En18 
    input [18:0] Wgt_0_58, // sfix19_En18 
    input [18:0] Wgt_0_59, // sfix19_En18 
    input [18:0] Wgt_0_60, // sfix19_En18 
    input [18:0] Wgt_0_61, // sfix19_En18 
    input [18:0] Wgt_0_62, // sfix19_En18 
    input [18:0] Wgt_0_63, // sfix19_En18 
    input [18:0] Wgt_0_64, // sfix19_En18 
    input [18:0] Wgt_0_65, // sfix19_En18 
    input [18:0] Wgt_0_66, // sfix19_En18 
    input [18:0] Wgt_0_67, // sfix19_En18 
    input [18:0] Wgt_0_68, // sfix19_En18 
    input [18:0] Wgt_0_69, // sfix19_En18 
    input [18:0] Wgt_0_70, // sfix19_En18 
    input [18:0] Wgt_0_71, // sfix19_En18 
    input [18:0] Wgt_0_72, // sfix19_En18 
    input [18:0] Wgt_0_73, // sfix19_En18 
    input [18:0] Wgt_0_74, // sfix19_En18 
    input [18:0] Wgt_0_75, // sfix19_En18 
    input [18:0] Wgt_0_76, // sfix19_En18 
    input [18:0] Wgt_0_77, // sfix19_En18 
    input [18:0] Wgt_0_78, // sfix19_En18 
    input [18:0] Wgt_0_79, // sfix19_En18 
    input [18:0] Wgt_0_80, // sfix19_En18 
    input [18:0] Wgt_0_81, // sfix19_En18 
    input [18:0] Wgt_0_82, // sfix19_En18 
    input [18:0] Wgt_0_83, // sfix19_En18 
    input [18:0] Wgt_0_84, // sfix19_En18 
    input [18:0] Wgt_0_85, // sfix19_En18 
    input [18:0] Wgt_0_86, // sfix19_En18 
    input [18:0] Wgt_0_87, // sfix19_En18 
    input [18:0] Wgt_0_88, // sfix19_En18 
    input [18:0] Wgt_0_89, // sfix19_En18 
    input [18:0] Wgt_0_90, // sfix19_En18 
    input [18:0] Wgt_0_91, // sfix19_En18 
    input [18:0] Wgt_0_92, // sfix19_En18 
    input [18:0] Wgt_0_93, // sfix19_En18 
    input [18:0] Wgt_0_94, // sfix19_En18 
    input [18:0] Wgt_0_95, // sfix19_En18 
    input [18:0] Wgt_0_96, // sfix19_En18 
    input [18:0] Wgt_0_97, // sfix19_En18 
    input [18:0] Wgt_0_98, // sfix19_En18 
    input [18:0] Wgt_0_99, // sfix19_En18 
    input [18:0] Wgt_0_100, // sfix19_En18 
    input [18:0] Wgt_0_101, // sfix19_En18 
    input [18:0] Wgt_0_102, // sfix19_En18 
    input [18:0] Wgt_0_103, // sfix19_En18 
    input [18:0] Wgt_0_104, // sfix19_En18 
    input [18:0] Wgt_0_105, // sfix19_En18 
    input [18:0] Wgt_0_106, // sfix19_En18 
    input [18:0] Wgt_0_107, // sfix19_En18 
    input [18:0] Wgt_0_108, // sfix19_En18 
    input [18:0] Wgt_0_109, // sfix19_En18 
    input [18:0] Wgt_0_110, // sfix19_En18 
    input [18:0] Wgt_0_111, // sfix19_En18 
    input [18:0] Wgt_0_112, // sfix19_En18 
    input [18:0] Wgt_0_113, // sfix19_En18 
    input [18:0] Wgt_0_114, // sfix19_En18 
    input [18:0] Wgt_0_115, // sfix19_En18 
    input [18:0] Wgt_0_116, // sfix19_En18 
    input [18:0] Wgt_0_117, // sfix19_En18 
    input [18:0] Wgt_0_118, // sfix19_En18 
    input [18:0] Wgt_0_119, // sfix19_En18 
    input [18:0] Wgt_0_120, // sfix19_En18 
    input [18:0] Wgt_0_121, // sfix19_En18 
    input [18:0] Wgt_0_122, // sfix19_En18 
    input [18:0] Wgt_0_123, // sfix19_En18 
    input [18:0] Wgt_0_124, // sfix19_En18 
    input [18:0] Wgt_0_125, // sfix19_En18 
    input [18:0] Wgt_0_126, // sfix19_En18 
    input [18:0] Wgt_0_127, // sfix19_En18 
    input [18:0] Wgt_0_128, // sfix19_En18 
    input [18:0] Wgt_0_129, // sfix19_En18 
    input [18:0] Wgt_0_130, // sfix19_En18 
    input [18:0] Wgt_0_131, // sfix19_En18 
    input [18:0] Wgt_0_132, // sfix19_En18 
    input [18:0] Wgt_0_133, // sfix19_En18 
    input [18:0] Wgt_0_134, // sfix19_En18 
    input [18:0] Wgt_0_135, // sfix19_En18 
    input [18:0] Wgt_0_136, // sfix19_En18 
    input [18:0] Wgt_0_137, // sfix19_En18 
    input [18:0] Wgt_0_138, // sfix19_En18 
    input [18:0] Wgt_0_139, // sfix19_En18 
    input [18:0] Wgt_0_140, // sfix19_En18 
    input [18:0] Wgt_0_141, // sfix19_En18 
    input [18:0] Wgt_0_142, // sfix19_En18 
    input [18:0] Wgt_0_143, // sfix19_En18 
    input [18:0] Wgt_0_144, // sfix19_En18 
    input [18:0] Wgt_0_145, // sfix19_En18 
    input [18:0] Wgt_0_146, // sfix19_En18 
    input [18:0] Wgt_0_147, // sfix19_En18 
    input [18:0] Wgt_0_148, // sfix19_En18 
    input [18:0] Wgt_0_149, // sfix19_En18 
    input [18:0] Wgt_0_150, // sfix19_En18 
    input [18:0] Wgt_0_151, // sfix19_En18 
    input [18:0] Wgt_0_152, // sfix19_En18 
    input [18:0] Wgt_0_153, // sfix19_En18 
    input [18:0] Wgt_0_154, // sfix19_En18 
    input [18:0] Wgt_0_155, // sfix19_En18 
    input [18:0] Wgt_0_156, // sfix19_En18 
    input [18:0] Wgt_0_157, // sfix19_En18 
    input [18:0] Wgt_0_158, // sfix19_En18 
    input [18:0] Wgt_0_159, // sfix19_En18 
    input [18:0] Wgt_0_160, // sfix19_En18 
    input [18:0] Wgt_0_161, // sfix19_En18 
    input [18:0] Wgt_0_162, // sfix19_En18 
    input [18:0] Wgt_0_163, // sfix19_En18 
    input [18:0] Wgt_0_164, // sfix19_En18 
    input [18:0] Wgt_0_165, // sfix19_En18 
    input [18:0] Wgt_0_166, // sfix19_En18 
    input [18:0] Wgt_0_167, // sfix19_En18 
    input [18:0] Wgt_0_168, // sfix19_En18 
    input [18:0] Wgt_0_169, // sfix19_En18 
    input [18:0] Wgt_0_170, // sfix19_En18 
    input [18:0] Wgt_0_171, // sfix19_En18 
    input [18:0] Wgt_0_172, // sfix19_En18 
    input [18:0] Wgt_0_173, // sfix19_En18 
    input [18:0] Wgt_0_174, // sfix19_En18 
    input [18:0] Wgt_0_175, // sfix19_En18 
    input [18:0] Wgt_0_176, // sfix19_En18 
    input [18:0] Wgt_0_177, // sfix19_En18 
    input [18:0] Wgt_0_178, // sfix19_En18 
    input [18:0] Wgt_0_179, // sfix19_En18 
    input [18:0] Wgt_0_180, // sfix19_En18 
    input [18:0] Wgt_0_181, // sfix19_En18 
    input [18:0] Wgt_0_182, // sfix19_En18 
    input [18:0] Wgt_0_183, // sfix19_En18 
    input [18:0] Wgt_0_184, // sfix19_En18 
    input [18:0] Wgt_0_185, // sfix19_En18 
    input [18:0] Wgt_0_186, // sfix19_En18 
    input [18:0] Wgt_0_187, // sfix19_En18 
    input [18:0] Wgt_0_188, // sfix19_En18 
    input [18:0] Wgt_0_189, // sfix19_En18 
    input [18:0] Wgt_0_190, // sfix19_En18 
    input [18:0] Wgt_0_191, // sfix19_En18 
    input [18:0] Wgt_0_192, // sfix19_En18 
    input [18:0] Wgt_0_193, // sfix19_En18 
    input [18:0] Wgt_0_194, // sfix19_En18 
    input [18:0] Wgt_0_195, // sfix19_En18 
    input [18:0] Wgt_0_196, // sfix19_En18 
    input [18:0] Wgt_0_197, // sfix19_En18 
    input [18:0] Wgt_0_198, // sfix19_En18 
    input [18:0] Wgt_0_199, // sfix19_En18 
    input [18:0] Wgt_0_200, // sfix19_En18 
    input [18:0] Wgt_0_201, // sfix19_En18 
    input [18:0] Wgt_0_202, // sfix19_En18 
    input [18:0] Wgt_0_203, // sfix19_En18 
    input [18:0] Wgt_0_204, // sfix19_En18 
    input [18:0] Wgt_0_205, // sfix19_En18 
    input [18:0] Wgt_0_206, // sfix19_En18 
    input [18:0] Wgt_0_207, // sfix19_En18 
    input [18:0] Wgt_0_208, // sfix19_En18 
    input [18:0] Wgt_0_209, // sfix19_En18 
    input [18:0] Wgt_0_210, // sfix19_En18 
    input [18:0] Wgt_0_211, // sfix19_En18 
    input [18:0] Wgt_0_212, // sfix19_En18 
    input [18:0] Wgt_0_213, // sfix19_En18 
    input [18:0] Wgt_0_214, // sfix19_En18 
    input [18:0] Wgt_0_215, // sfix19_En18 
    input [18:0] Wgt_0_216, // sfix19_En18 
    input [18:0] Wgt_0_217, // sfix19_En18 
    input [18:0] Wgt_0_218, // sfix19_En18 
    input [18:0] Wgt_0_219, // sfix19_En18 
    input [18:0] Wgt_0_220, // sfix19_En18 
    input [18:0] Wgt_0_221, // sfix19_En18 
    input [18:0] Wgt_0_222, // sfix19_En18 
    input [18:0] Wgt_0_223, // sfix19_En18 
    input [18:0] Wgt_0_224, // sfix19_En18 
    input [18:0] Wgt_0_225, // sfix19_En18 
    input [18:0] Wgt_0_226, // sfix19_En18 
    input [18:0] Wgt_0_227, // sfix19_En18 
    input [18:0] Wgt_0_228, // sfix19_En18 
    input [18:0] Wgt_0_229, // sfix19_En18 
    input [18:0] Wgt_0_230, // sfix19_En18 
    input [18:0] Wgt_0_231, // sfix19_En18 
    input [18:0] Wgt_0_232, // sfix19_En18 
    input [18:0] Wgt_0_233, // sfix19_En18 
    input [18:0] Wgt_0_234, // sfix19_En18 
    input [18:0] Wgt_0_235, // sfix19_En18 
    input [18:0] Wgt_0_236, // sfix19_En18 
    input [18:0] Wgt_0_237, // sfix19_En18 
    input [18:0] Wgt_0_238, // sfix19_En18 
    input [18:0] Wgt_0_239, // sfix19_En18 
    input [18:0] Wgt_0_240, // sfix19_En18 
    input [18:0] Wgt_0_241, // sfix19_En18 
    input [18:0] Wgt_0_242, // sfix19_En18 
    input [18:0] Wgt_0_243, // sfix19_En18 
    input [18:0] Wgt_0_244, // sfix19_En18 
    input [18:0] Wgt_0_245, // sfix19_En18 
    input [18:0] Wgt_0_246, // sfix19_En18 
    input [18:0] Wgt_0_247, // sfix19_En18 
    input [18:0] Wgt_0_248, // sfix19_En18 
    input [18:0] Wgt_0_249, // sfix19_En18 
    input [18:0] Wgt_0_250, // sfix19_En18 
    input [18:0] Wgt_0_251, // sfix19_En18 
    input [18:0] Wgt_0_252, // sfix19_En18 
    input [18:0] Wgt_0_253, // sfix19_En18 
    input [18:0] Wgt_0_254, // sfix19_En18 
    input [18:0] Wgt_0_255, // sfix19_En18 
    input [18:0] Wgt_0_256, // sfix19_En18 
    input [18:0] Wgt_0_257, // sfix19_En18 
    input [18:0] Wgt_0_258, // sfix19_En18 
    input [18:0] Wgt_0_259, // sfix19_En18 
    input [18:0] Wgt_0_260, // sfix19_En18 
    input [18:0] Wgt_0_261, // sfix19_En18 
    input [18:0] Wgt_0_262, // sfix19_En18 
    input [18:0] Wgt_0_263, // sfix19_En18 
    input [18:0] Wgt_0_264, // sfix19_En18 
    input [18:0] Wgt_0_265, // sfix19_En18 
    input [18:0] Wgt_0_266, // sfix19_En18 
    input [18:0] Wgt_0_267, // sfix19_En18 
    input [18:0] Wgt_0_268, // sfix19_En18 
    input [18:0] Wgt_0_269, // sfix19_En18 
    input [18:0] Wgt_0_270, // sfix19_En18 
    input [18:0] Wgt_0_271, // sfix19_En18 
    input [18:0] Wgt_0_272, // sfix19_En18 
    input [18:0] Wgt_0_273, // sfix19_En18 
    input [18:0] Wgt_0_274, // sfix19_En18 
    input [18:0] Wgt_0_275, // sfix19_En18 
    input [18:0] Wgt_0_276, // sfix19_En18 
    input [18:0] Wgt_0_277, // sfix19_En18 
    input [18:0] Wgt_0_278, // sfix19_En18 
    input [18:0] Wgt_0_279, // sfix19_En18 
    input [18:0] Wgt_0_280, // sfix19_En18 
    input [18:0] Wgt_0_281, // sfix19_En18 
    input [18:0] Wgt_0_282, // sfix19_En18 
    input [18:0] Wgt_0_283, // sfix19_En18 
    input [18:0] Wgt_0_284, // sfix19_En18 
    input [18:0] Wgt_0_285, // sfix19_En18 
    input [18:0] Wgt_0_286, // sfix19_En18 
    input [18:0] Wgt_0_287, // sfix19_En18 
    input [18:0] Wgt_0_288, // sfix19_En18 
    input [18:0] Wgt_0_289, // sfix19_En18 
    input [18:0] Wgt_0_290, // sfix19_En18 
    input [18:0] Wgt_0_291, // sfix19_En18 
    input [18:0] Wgt_0_292, // sfix19_En18 
    input [18:0] Wgt_0_293, // sfix19_En18 
    input [18:0] Wgt_0_294, // sfix19_En18 
    input [18:0] Wgt_0_295, // sfix19_En18 
    input [18:0] Wgt_0_296, // sfix19_En18 
    input [18:0] Wgt_0_297, // sfix19_En18 
    input [18:0] Wgt_0_298, // sfix19_En18 
    input [18:0] Wgt_0_299, // sfix19_En18 
    input [18:0] Wgt_0_300, // sfix19_En18 
    input [18:0] Wgt_0_301, // sfix19_En18 
    input [18:0] Wgt_0_302, // sfix19_En18 
    input [18:0] Wgt_0_303, // sfix19_En18 
    input [18:0] Wgt_0_304, // sfix19_En18 
    input [18:0] Wgt_0_305, // sfix19_En18 
    input [18:0] Wgt_0_306, // sfix19_En18 
    input [18:0] Wgt_0_307, // sfix19_En18 
    input [18:0] Wgt_0_308, // sfix19_En18 
    input [18:0] Wgt_0_309, // sfix19_En18 
    input [18:0] Wgt_0_310, // sfix19_En18 
    input [18:0] Wgt_0_311, // sfix19_En18 
    input [18:0] Wgt_0_312, // sfix19_En18 
    input [18:0] Wgt_0_313, // sfix19_En18 
    input [18:0] Wgt_0_314, // sfix19_En18 
    input [18:0] Wgt_0_315, // sfix19_En18 
    input [18:0] Wgt_0_316, // sfix19_En18 
    input [18:0] Wgt_0_317, // sfix19_En18 
    input [18:0] Wgt_0_318, // sfix19_En18 
    input [18:0] Wgt_0_319, // sfix19_En18 
    input [18:0] Wgt_0_320, // sfix19_En18 
    input [18:0] Wgt_0_321, // sfix19_En18 
    input [18:0] Wgt_0_322, // sfix19_En18 
    input [18:0] Wgt_0_323, // sfix19_En18 
    input [18:0] Wgt_0_324, // sfix19_En18 
    input [18:0] Wgt_0_325, // sfix19_En18 
    input [18:0] Wgt_0_326, // sfix19_En18 
    input [18:0] Wgt_0_327, // sfix19_En18 
    input [18:0] Wgt_0_328, // sfix19_En18 
    input [18:0] Wgt_0_329, // sfix19_En18 
    input [18:0] Wgt_0_330, // sfix19_En18 
    input [18:0] Wgt_0_331, // sfix19_En18 
    input [18:0] Wgt_0_332, // sfix19_En18 
    input [18:0] Wgt_0_333, // sfix19_En18 
    input [18:0] Wgt_0_334, // sfix19_En18 
    input [18:0] Wgt_0_335, // sfix19_En18 
    input [18:0] Wgt_0_336, // sfix19_En18 
    input [18:0] Wgt_0_337, // sfix19_En18 
    input [18:0] Wgt_0_338, // sfix19_En18 
    input [18:0] Wgt_0_339, // sfix19_En18 
    input [18:0] Wgt_0_340, // sfix19_En18 
    input [18:0] Wgt_0_341, // sfix19_En18 
    input [18:0] Wgt_0_342, // sfix19_En18 
    input [18:0] Wgt_0_343, // sfix19_En18 
    input [18:0] Wgt_0_344, // sfix19_En18 
    input [18:0] Wgt_0_345, // sfix19_En18 
    input [18:0] Wgt_0_346, // sfix19_En18 
    input [18:0] Wgt_0_347, // sfix19_En18 
    input [18:0] Wgt_0_348, // sfix19_En18 
    input [18:0] Wgt_0_349, // sfix19_En18 
    input [18:0] Wgt_0_350, // sfix19_En18 
    input [18:0] Wgt_0_351, // sfix19_En18 
    input [18:0] Wgt_0_352, // sfix19_En18 
    input [18:0] Wgt_0_353, // sfix19_En18 
    input [18:0] Wgt_0_354, // sfix19_En18 
    input [18:0] Wgt_0_355, // sfix19_En18 
    input [18:0] Wgt_0_356, // sfix19_En18 
    input [18:0] Wgt_0_357, // sfix19_En18 
    input [18:0] Wgt_0_358, // sfix19_En18 
    input [18:0] Wgt_0_359, // sfix19_En18 
    input [18:0] Wgt_0_360, // sfix19_En18 
    input [18:0] Wgt_0_361, // sfix19_En18 
    input [18:0] Wgt_0_362, // sfix19_En18 
    input [18:0] Wgt_0_363, // sfix19_En18 
    input [18:0] Wgt_0_364, // sfix19_En18 
    input [18:0] Wgt_0_365, // sfix19_En18 
    input [18:0] Wgt_0_366, // sfix19_En18 
    input [18:0] Wgt_0_367, // sfix19_En18 
    input [18:0] Wgt_0_368, // sfix19_En18 
    input [18:0] Wgt_0_369, // sfix19_En18 
    input [18:0] Wgt_0_370, // sfix19_En18 
    input [18:0] Wgt_0_371, // sfix19_En18 
    input [18:0] Wgt_0_372, // sfix19_En18 
    input [18:0] Wgt_0_373, // sfix19_En18 
    input [18:0] Wgt_0_374, // sfix19_En18 
    input [18:0] Wgt_0_375, // sfix19_En18 
    input [18:0] Wgt_0_376, // sfix19_En18 
    input [18:0] Wgt_0_377, // sfix19_En18 
    input [18:0] Wgt_0_378, // sfix19_En18 
    input [18:0] Wgt_0_379, // sfix19_En18 
    input [18:0] Wgt_0_380, // sfix19_En18 
    input [18:0] Wgt_0_381, // sfix19_En18 
    input [18:0] Wgt_0_382, // sfix19_En18 
    input [18:0] Wgt_0_383, // sfix19_En18 
    input [18:0] Wgt_0_384, // sfix19_En18 
    input [18:0] Wgt_0_385, // sfix19_En18 
    input [18:0] Wgt_0_386, // sfix19_En18 
    input [18:0] Wgt_0_387, // sfix19_En18 
    input [18:0] Wgt_0_388, // sfix19_En18 
    input [18:0] Wgt_0_389, // sfix19_En18 
    input [18:0] Wgt_0_390, // sfix19_En18 
    input [18:0] Wgt_0_391, // sfix19_En18 
    input [18:0] Wgt_0_392, // sfix19_En18 
    input [18:0] Wgt_0_393, // sfix19_En18 
    input [18:0] Wgt_0_394, // sfix19_En18 
    input [18:0] Wgt_0_395, // sfix19_En18 
    input [18:0] Wgt_0_396, // sfix19_En18 
    input [18:0] Wgt_0_397, // sfix19_En18 
    input [18:0] Wgt_0_398, // sfix19_En18 
    input [18:0] Wgt_0_399, // sfix19_En18 
    input [18:0] Wgt_0_400, // sfix19_En18 
    input [18:0] Wgt_0_401, // sfix19_En18 
    input [18:0] Wgt_0_402, // sfix19_En18 
    input [18:0] Wgt_0_403, // sfix19_En18 
    input [18:0] Wgt_0_404, // sfix19_En18 
    input [18:0] Wgt_0_405, // sfix19_En18 
    input [18:0] Wgt_0_406, // sfix19_En18 
    input [18:0] Wgt_0_407, // sfix19_En18 
    input [18:0] Wgt_0_408, // sfix19_En18 
    input [18:0] Wgt_0_409, // sfix19_En18 
    input [18:0] Wgt_0_410, // sfix19_En18 
    input [18:0] Wgt_0_411, // sfix19_En18 
    input [18:0] Wgt_0_412, // sfix19_En18 
    input [18:0] Wgt_0_413, // sfix19_En18 
    input [18:0] Wgt_0_414, // sfix19_En18 
    input [18:0] Wgt_0_415, // sfix19_En18 
    input [18:0] Wgt_0_416, // sfix19_En18 
    input [18:0] Wgt_0_417, // sfix19_En18 
    input [18:0] Wgt_0_418, // sfix19_En18 
    input [18:0] Wgt_0_419, // sfix19_En18 
    input [18:0] Wgt_0_420, // sfix19_En18 
    input [18:0] Wgt_0_421, // sfix19_En18 
    input [18:0] Wgt_0_422, // sfix19_En18 
    input [18:0] Wgt_0_423, // sfix19_En18 
    input [18:0] Wgt_0_424, // sfix19_En18 
    input [18:0] Wgt_0_425, // sfix19_En18 
    input [18:0] Wgt_0_426, // sfix19_En18 
    input [18:0] Wgt_0_427, // sfix19_En18 
    input [18:0] Wgt_0_428, // sfix19_En18 
    input [18:0] Wgt_0_429, // sfix19_En18 
    input [18:0] Wgt_0_430, // sfix19_En18 
    input [18:0] Wgt_0_431, // sfix19_En18 
    input [18:0] Wgt_0_432, // sfix19_En18 
    input [18:0] Wgt_0_433, // sfix19_En18 
    input [18:0] Wgt_0_434, // sfix19_En18 
    input [18:0] Wgt_0_435, // sfix19_En18 
    input [18:0] Wgt_0_436, // sfix19_En18 
    input [18:0] Wgt_0_437, // sfix19_En18 
    input [18:0] Wgt_0_438, // sfix19_En18 
    input [18:0] Wgt_0_439, // sfix19_En18 
    input [18:0] Wgt_0_440, // sfix19_En18 
    input [18:0] Wgt_0_441, // sfix19_En18 
    input [18:0] Wgt_0_442, // sfix19_En18 
    input [18:0] Wgt_0_443, // sfix19_En18 
    input [18:0] Wgt_0_444, // sfix19_En18 
    input [18:0] Wgt_0_445, // sfix19_En18 
    input [18:0] Wgt_0_446, // sfix19_En18 
    input [18:0] Wgt_0_447, // sfix19_En18 
    input [18:0] Wgt_0_448, // sfix19_En18 
    input [18:0] Wgt_0_449, // sfix19_En18 
    input [18:0] Wgt_0_450, // sfix19_En18 
    input [18:0] Wgt_0_451, // sfix19_En18 
    input [18:0] Wgt_0_452, // sfix19_En18 
    input [18:0] Wgt_0_453, // sfix19_En18 
    input [18:0] Wgt_0_454, // sfix19_En18 
    input [18:0] Wgt_0_455, // sfix19_En18 
    input [18:0] Wgt_0_456, // sfix19_En18 
    input [18:0] Wgt_0_457, // sfix19_En18 
    input [18:0] Wgt_0_458, // sfix19_En18 
    input [18:0] Wgt_0_459, // sfix19_En18 
    input [18:0] Wgt_0_460, // sfix19_En18 
    input [18:0] Wgt_0_461, // sfix19_En18 
    input [18:0] Wgt_0_462, // sfix19_En18 
    input [18:0] Wgt_0_463, // sfix19_En18 
    input [18:0] Wgt_0_464, // sfix19_En18 
    input [18:0] Wgt_0_465, // sfix19_En18 
    input [18:0] Wgt_0_466, // sfix19_En18 
    input [18:0] Wgt_0_467, // sfix19_En18 
    input [18:0] Wgt_0_468, // sfix19_En18 
    input [18:0] Wgt_0_469, // sfix19_En18 
    input [18:0] Wgt_0_470, // sfix19_En18 
    input [18:0] Wgt_0_471, // sfix19_En18 
    input [18:0] Wgt_0_472, // sfix19_En18 
    input [18:0] Wgt_0_473, // sfix19_En18 
    input [18:0] Wgt_0_474, // sfix19_En18 
    input [18:0] Wgt_0_475, // sfix19_En18 
    input [18:0] Wgt_0_476, // sfix19_En18 
    input [18:0] Wgt_0_477, // sfix19_En18 
    input [18:0] Wgt_0_478, // sfix19_En18 
    input [18:0] Wgt_0_479, // sfix19_En18 
    input [18:0] Wgt_0_480, // sfix19_En18 
    input [18:0] Wgt_0_481, // sfix19_En18 
    input [18:0] Wgt_0_482, // sfix19_En18 
    input [18:0] Wgt_0_483, // sfix19_En18 
    input [18:0] Wgt_0_484, // sfix19_En18 
    input [18:0] Wgt_0_485, // sfix19_En18 
    input [18:0] Wgt_0_486, // sfix19_En18 
    input [18:0] Wgt_0_487, // sfix19_En18 
    input [18:0] Wgt_0_488, // sfix19_En18 
    input [18:0] Wgt_0_489, // sfix19_En18 
    input [18:0] Wgt_0_490, // sfix19_En18 
    input [18:0] Wgt_0_491, // sfix19_En18 
    input [18:0] Wgt_0_492, // sfix19_En18 
    input [18:0] Wgt_0_493, // sfix19_En18 
    input [18:0] Wgt_0_494, // sfix19_En18 
    input [18:0] Wgt_0_495, // sfix19_En18 
    input [18:0] Wgt_0_496, // sfix19_En18 
    input [18:0] Wgt_0_497, // sfix19_En18 
    input [18:0] Wgt_0_498, // sfix19_En18 
    input [18:0] Wgt_0_499, // sfix19_En18 
    input [18:0] Wgt_0_500, // sfix19_En18 
    input [18:0] Wgt_0_501, // sfix19_En18 
    input [18:0] Wgt_0_502, // sfix19_En18 
    input [18:0] Wgt_0_503, // sfix19_En18 
    input [18:0] Wgt_0_504, // sfix19_En18 
    input [18:0] Wgt_0_505, // sfix19_En18 
    input [18:0] Wgt_0_506, // sfix19_En18 
    input [18:0] Wgt_0_507, // sfix19_En18 
    input [18:0] Wgt_0_508, // sfix19_En18 
    input [18:0] Wgt_0_509, // sfix19_En18 
    input [18:0] Wgt_0_510, // sfix19_En18 
    input [18:0] Wgt_0_511, // sfix19_En18 
    input [18:0] Wgt_0_512, // sfix19_En18 
    input [18:0] Wgt_0_513, // sfix19_En18 
    input [18:0] Wgt_0_514, // sfix19_En18 
    input [18:0] Wgt_0_515, // sfix19_En18 
    input [18:0] Wgt_0_516, // sfix19_En18 
    input [18:0] Wgt_0_517, // sfix19_En18 
    input [18:0] Wgt_0_518, // sfix19_En18 
    input [18:0] Wgt_0_519, // sfix19_En18 
    input [18:0] Wgt_0_520, // sfix19_En18 
    input [18:0] Wgt_0_521, // sfix19_En18 
    input [18:0] Wgt_0_522, // sfix19_En18 
    input [18:0] Wgt_0_523, // sfix19_En18 
    input [18:0] Wgt_0_524, // sfix19_En18 
    input [18:0] Wgt_0_525, // sfix19_En18 
    input [18:0] Wgt_0_526, // sfix19_En18 
    input [18:0] Wgt_0_527, // sfix19_En18 
    input [18:0] Wgt_0_528, // sfix19_En18 
    input [18:0] Wgt_0_529, // sfix19_En18 
    input [18:0] Wgt_0_530, // sfix19_En18 
    input [18:0] Wgt_0_531, // sfix19_En18 
    input [18:0] Wgt_0_532, // sfix19_En18 
    input [18:0] Wgt_0_533, // sfix19_En18 
    input [18:0] Wgt_0_534, // sfix19_En18 
    input [18:0] Wgt_0_535, // sfix19_En18 
    input [18:0] Wgt_0_536, // sfix19_En18 
    input [18:0] Wgt_0_537, // sfix19_En18 
    input [18:0] Wgt_0_538, // sfix19_En18 
    input [18:0] Wgt_0_539, // sfix19_En18 
    input [18:0] Wgt_0_540, // sfix19_En18 
    input [18:0] Wgt_0_541, // sfix19_En18 
    input [18:0] Wgt_0_542, // sfix19_En18 
    input [18:0] Wgt_0_543, // sfix19_En18 
    input [18:0] Wgt_0_544, // sfix19_En18 
    input [18:0] Wgt_0_545, // sfix19_En18 
    input [18:0] Wgt_0_546, // sfix19_En18 
    input [18:0] Wgt_0_547, // sfix19_En18 
    input [18:0] Wgt_0_548, // sfix19_En18 
    input [18:0] Wgt_0_549, // sfix19_En18 
    input [18:0] Wgt_0_550, // sfix19_En18 
    input [18:0] Wgt_0_551, // sfix19_En18 
    input [18:0] Wgt_0_552, // sfix19_En18 
    input [18:0] Wgt_0_553, // sfix19_En18 
    input [18:0] Wgt_0_554, // sfix19_En18 
    input [18:0] Wgt_0_555, // sfix19_En18 
    input [18:0] Wgt_0_556, // sfix19_En18 
    input [18:0] Wgt_0_557, // sfix19_En18 
    input [18:0] Wgt_0_558, // sfix19_En18 
    input [18:0] Wgt_0_559, // sfix19_En18 
    input [18:0] Wgt_0_560, // sfix19_En18 
    input [18:0] Wgt_0_561, // sfix19_En18 
    input [18:0] Wgt_0_562, // sfix19_En18 
    input [18:0] Wgt_0_563, // sfix19_En18 
    input [18:0] Wgt_0_564, // sfix19_En18 
    input [18:0] Wgt_0_565, // sfix19_En18 
    input [18:0] Wgt_0_566, // sfix19_En18 
    input [18:0] Wgt_0_567, // sfix19_En18 
    input [18:0] Wgt_0_568, // sfix19_En18 
    input [18:0] Wgt_0_569, // sfix19_En18 
    input [18:0] Wgt_0_570, // sfix19_En18 
    input [18:0] Wgt_0_571, // sfix19_En18 
    input [18:0] Wgt_0_572, // sfix19_En18 
    input [18:0] Wgt_0_573, // sfix19_En18 
    input [18:0] Wgt_0_574, // sfix19_En18 
    input [18:0] Wgt_0_575, // sfix19_En18 
    input [18:0] Wgt_0_576, // sfix19_En18 
    input [18:0] Wgt_0_577, // sfix19_En18 
    input [18:0] Wgt_0_578, // sfix19_En18 
    input [18:0] Wgt_0_579, // sfix19_En18 
    input [18:0] Wgt_0_580, // sfix19_En18 
    input [18:0] Wgt_0_581, // sfix19_En18 
    input [18:0] Wgt_0_582, // sfix19_En18 
    input [18:0] Wgt_0_583, // sfix19_En18 
    input [18:0] Wgt_0_584, // sfix19_En18 
    input [18:0] Wgt_0_585, // sfix19_En18 
    input [18:0] Wgt_0_586, // sfix19_En18 
    input [18:0] Wgt_0_587, // sfix19_En18 
    input [18:0] Wgt_0_588, // sfix19_En18 
    input [18:0] Wgt_0_589, // sfix19_En18 
    input [18:0] Wgt_0_590, // sfix19_En18 
    input [18:0] Wgt_0_591, // sfix19_En18 
    input [18:0] Wgt_0_592, // sfix19_En18 
    input [18:0] Wgt_0_593, // sfix19_En18 
    input [18:0] Wgt_0_594, // sfix19_En18 
    input [18:0] Wgt_0_595, // sfix19_En18 
    input [18:0] Wgt_0_596, // sfix19_En18 
    input [18:0] Wgt_0_597, // sfix19_En18 
    input [18:0] Wgt_0_598, // sfix19_En18 
    input [18:0] Wgt_0_599, // sfix19_En18 
    input [18:0] Wgt_0_600, // sfix19_En18 
    input [18:0] Wgt_0_601, // sfix19_En18 
    input [18:0] Wgt_0_602, // sfix19_En18 
    input [18:0] Wgt_0_603, // sfix19_En18 
    input [18:0] Wgt_0_604, // sfix19_En18 
    input [18:0] Wgt_0_605, // sfix19_En18 
    input [18:0] Wgt_0_606, // sfix19_En18 
    input [18:0] Wgt_0_607, // sfix19_En18 
    input [18:0] Wgt_0_608, // sfix19_En18 
    input [18:0] Wgt_0_609, // sfix19_En18 
    input [18:0] Wgt_0_610, // sfix19_En18 
    input [18:0] Wgt_0_611, // sfix19_En18 
    input [18:0] Wgt_0_612, // sfix19_En18 
    input [18:0] Wgt_0_613, // sfix19_En18 
    input [18:0] Wgt_0_614, // sfix19_En18 
    input [18:0] Wgt_0_615, // sfix19_En18 
    input [18:0] Wgt_0_616, // sfix19_En18 
    input [18:0] Wgt_0_617, // sfix19_En18 
    input [18:0] Wgt_0_618, // sfix19_En18 
    input [18:0] Wgt_0_619, // sfix19_En18 
    input [18:0] Wgt_0_620, // sfix19_En18 
    input [18:0] Wgt_0_621, // sfix19_En18 
    input [18:0] Wgt_0_622, // sfix19_En18 
    input [18:0] Wgt_0_623, // sfix19_En18 
    input [18:0] Wgt_0_624, // sfix19_En18 
    input [18:0] Wgt_0_625, // sfix19_En18 
    input [18:0] Wgt_0_626, // sfix19_En18 
    input [18:0] Wgt_0_627, // sfix19_En18 
    input [18:0] Wgt_0_628, // sfix19_En18 
    input [18:0] Wgt_0_629, // sfix19_En18 
    input [18:0] Wgt_0_630, // sfix19_En18 
    input [18:0] Wgt_0_631, // sfix19_En18 
    input [18:0] Wgt_0_632, // sfix19_En18 
    input [18:0] Wgt_0_633, // sfix19_En18 
    input [18:0] Wgt_0_634, // sfix19_En18 
    input [18:0] Wgt_0_635, // sfix19_En18 
    input [18:0] Wgt_0_636, // sfix19_En18 
    input [18:0] Wgt_0_637, // sfix19_En18 
    input [18:0] Wgt_0_638, // sfix19_En18 
    input [18:0] Wgt_0_639, // sfix19_En18 
    input [18:0] Wgt_0_640, // sfix19_En18 
    input [18:0] Wgt_0_641, // sfix19_En18 
    input [18:0] Wgt_0_642, // sfix19_En18 
    input [18:0] Wgt_0_643, // sfix19_En18 
    input [18:0] Wgt_0_644, // sfix19_En18 
    input [18:0] Wgt_0_645, // sfix19_En18 
    input [18:0] Wgt_0_646, // sfix19_En18 
    input [18:0] Wgt_0_647, // sfix19_En18 
    input [18:0] Wgt_0_648, // sfix19_En18 
    input [18:0] Wgt_0_649, // sfix19_En18 
    input [18:0] Wgt_0_650, // sfix19_En18 
    input [18:0] Wgt_0_651, // sfix19_En18 
    input [18:0] Wgt_0_652, // sfix19_En18 
    input [18:0] Wgt_0_653, // sfix19_En18 
    input [18:0] Wgt_0_654, // sfix19_En18 
    input [18:0] Wgt_0_655, // sfix19_En18 
    input [18:0] Wgt_0_656, // sfix19_En18 
    input [18:0] Wgt_0_657, // sfix19_En18 
    input [18:0] Wgt_0_658, // sfix19_En18 
    input [18:0] Wgt_0_659, // sfix19_En18 
    input [18:0] Wgt_0_660, // sfix19_En18 
    input [18:0] Wgt_0_661, // sfix19_En18 
    input [18:0] Wgt_0_662, // sfix19_En18 
    input [18:0] Wgt_0_663, // sfix19_En18 
    input [18:0] Wgt_0_664, // sfix19_En18 
    input [18:0] Wgt_0_665, // sfix19_En18 
    input [18:0] Wgt_0_666, // sfix19_En18 
    input [18:0] Wgt_0_667, // sfix19_En18 
    input [18:0] Wgt_0_668, // sfix19_En18 
    input [18:0] Wgt_0_669, // sfix19_En18 
    input [18:0] Wgt_0_670, // sfix19_En18 
    input [18:0] Wgt_0_671, // sfix19_En18 
    input [18:0] Wgt_0_672, // sfix19_En18 
    input [18:0] Wgt_0_673, // sfix19_En18 
    input [18:0] Wgt_0_674, // sfix19_En18 
    input [18:0] Wgt_0_675, // sfix19_En18 
    input [18:0] Wgt_0_676, // sfix19_En18 
    input [18:0] Wgt_0_677, // sfix19_En18 
    input [18:0] Wgt_0_678, // sfix19_En18 
    input [18:0] Wgt_0_679, // sfix19_En18 
    input [18:0] Wgt_0_680, // sfix19_En18 
    input [18:0] Wgt_0_681, // sfix19_En18 
    input [18:0] Wgt_0_682, // sfix19_En18 
    input [18:0] Wgt_0_683, // sfix19_En18 
    input [18:0] Wgt_0_684, // sfix19_En18 
    input [18:0] Wgt_0_685, // sfix19_En18 
    input [18:0] Wgt_0_686, // sfix19_En18 
    input [18:0] Wgt_0_687, // sfix19_En18 
    input [18:0] Wgt_0_688, // sfix19_En18 
    input [18:0] Wgt_0_689, // sfix19_En18 
    input [18:0] Wgt_0_690, // sfix19_En18 
    input [18:0] Wgt_0_691, // sfix19_En18 
    input [18:0] Wgt_0_692, // sfix19_En18 
    input [18:0] Wgt_0_693, // sfix19_En18 
    input [18:0] Wgt_0_694, // sfix19_En18 
    input [18:0] Wgt_0_695, // sfix19_En18 
    input [18:0] Wgt_0_696, // sfix19_En18 
    input [18:0] Wgt_0_697, // sfix19_En18 
    input [18:0] Wgt_0_698, // sfix19_En18 
    input [18:0] Wgt_0_699, // sfix19_En18 
    input [18:0] Wgt_0_700, // sfix19_En18 
    input [18:0] Wgt_0_701, // sfix19_En18 
    input [18:0] Wgt_0_702, // sfix19_En18 
    input [18:0] Wgt_0_703, // sfix19_En18 
    input [18:0] Wgt_0_704, // sfix19_En18 
    input [18:0] Wgt_0_705, // sfix19_En18 
    input [18:0] Wgt_0_706, // sfix19_En18 
    input [18:0] Wgt_0_707, // sfix19_En18 
    input [18:0] Wgt_0_708, // sfix19_En18 
    input [18:0] Wgt_0_709, // sfix19_En18 
    input [18:0] Wgt_0_710, // sfix19_En18 
    input [18:0] Wgt_0_711, // sfix19_En18 
    input [18:0] Wgt_0_712, // sfix19_En18 
    input [18:0] Wgt_0_713, // sfix19_En18 
    input [18:0] Wgt_0_714, // sfix19_En18 
    input [18:0] Wgt_0_715, // sfix19_En18 
    input [18:0] Wgt_0_716, // sfix19_En18 
    input [18:0] Wgt_0_717, // sfix19_En18 
    input [18:0] Wgt_0_718, // sfix19_En18 
    input [18:0] Wgt_0_719, // sfix19_En18 
    input [18:0] Wgt_0_720, // sfix19_En18 
    input [18:0] Wgt_0_721, // sfix19_En18 
    input [18:0] Wgt_0_722, // sfix19_En18 
    input [18:0] Wgt_0_723, // sfix19_En18 
    input [18:0] Wgt_0_724, // sfix19_En18 
    input [18:0] Wgt_0_725, // sfix19_En18 
    input [18:0] Wgt_0_726, // sfix19_En18 
    input [18:0] Wgt_0_727, // sfix19_En18 
    input [18:0] Wgt_0_728, // sfix19_En18 
    input [18:0] Wgt_0_729, // sfix19_En18 
    input [18:0] Wgt_0_730, // sfix19_En18 
    input [18:0] Wgt_0_731, // sfix19_En18 
    input [18:0] Wgt_0_732, // sfix19_En18 
    input [18:0] Wgt_0_733, // sfix19_En18 
    input [18:0] Wgt_0_734, // sfix19_En18 
    input [18:0] Wgt_0_735, // sfix19_En18 
    input [18:0] Wgt_0_736, // sfix19_En18 
    input [18:0] Wgt_0_737, // sfix19_En18 
    input [18:0] Wgt_0_738, // sfix19_En18 
    input [18:0] Wgt_0_739, // sfix19_En18 
    input [18:0] Wgt_0_740, // sfix19_En18 
    input [18:0] Wgt_0_741, // sfix19_En18 
    input [18:0] Wgt_0_742, // sfix19_En18 
    input [18:0] Wgt_0_743, // sfix19_En18 
    input [18:0] Wgt_0_744, // sfix19_En18 
    input [18:0] Wgt_0_745, // sfix19_En18 
    input [18:0] Wgt_0_746, // sfix19_En18 
    input [18:0] Wgt_0_747, // sfix19_En18 
    input [18:0] Wgt_0_748, // sfix19_En18 
    input [18:0] Wgt_0_749, // sfix19_En18 
    input [18:0] Wgt_0_750, // sfix19_En18 
    input [18:0] Wgt_0_751, // sfix19_En18 
    input [18:0] Wgt_0_752, // sfix19_En18 
    input [18:0] Wgt_0_753, // sfix19_En18 
    input [18:0] Wgt_0_754, // sfix19_En18 
    input [18:0] Wgt_0_755, // sfix19_En18 
    input [18:0] Wgt_0_756, // sfix19_En18 
    input [18:0] Wgt_0_757, // sfix19_En18 
    input [18:0] Wgt_0_758, // sfix19_En18 
    input [18:0] Wgt_0_759, // sfix19_En18 
    input [18:0] Wgt_0_760, // sfix19_En18 
    input [18:0] Wgt_0_761, // sfix19_En18 
    input [18:0] Wgt_0_762, // sfix19_En18 
    input [18:0] Wgt_0_763, // sfix19_En18 
    input [18:0] Wgt_0_764, // sfix19_En18 
    input [18:0] Wgt_0_765, // sfix19_En18 
    input [18:0] Wgt_0_766, // sfix19_En18 
    input [18:0] Wgt_0_767, // sfix19_En18 
    input [18:0] Wgt_0_768, // sfix19_En18 
    input [18:0] Wgt_0_769, // sfix19_En18 
    input [18:0] Wgt_0_770, // sfix19_En18 
    input [18:0] Wgt_0_771, // sfix19_En18 
    input [18:0] Wgt_0_772, // sfix19_En18 
    input [18:0] Wgt_0_773, // sfix19_En18 
    input [18:0] Wgt_0_774, // sfix19_En18 
    input [18:0] Wgt_0_775, // sfix19_En18 
    input [18:0] Wgt_0_776, // sfix19_En18 
    input [18:0] Wgt_0_777, // sfix19_En18 
    input [18:0] Wgt_0_778, // sfix19_En18 
    input [18:0] Wgt_0_779, // sfix19_En18 
    input [18:0] Wgt_0_780, // sfix19_En18 
    input [18:0] Wgt_0_781, // sfix19_En18 
    input [18:0] Wgt_0_782, // sfix19_En18 
    input [18:0] Wgt_0_783, // sfix19_En18 
    input [18:0] Wgt_0_784, // sfix19_En18 
    input [18:0] Wgt_1_0, // sfix19_En18 
    input [18:0] Wgt_1_1, // sfix19_En18 
    input [18:0] Wgt_1_2, // sfix19_En18 
    input [18:0] Wgt_1_3, // sfix19_En18 
    input [18:0] Wgt_1_4, // sfix19_En18 
    input [18:0] Wgt_1_5, // sfix19_En18 
    input [18:0] Wgt_1_6, // sfix19_En18 
    input [18:0] Wgt_1_7, // sfix19_En18 
    input [18:0] Wgt_1_8, // sfix19_En18 
    input [18:0] Wgt_1_9, // sfix19_En18 
    input [18:0] Wgt_1_10, // sfix19_En18 
    input [18:0] Wgt_1_11, // sfix19_En18 
    input [18:0] Wgt_1_12, // sfix19_En18 
    input [18:0] Wgt_1_13, // sfix19_En18 
    input [18:0] Wgt_1_14, // sfix19_En18 
    input [18:0] Wgt_1_15, // sfix19_En18 
    input [18:0] Wgt_1_16, // sfix19_En18 
    input [18:0] Wgt_1_17, // sfix19_En18 
    input [18:0] Wgt_1_18, // sfix19_En18 
    input [18:0] Wgt_1_19, // sfix19_En18 
    input [18:0] Wgt_1_20, // sfix19_En18 
    input [18:0] Wgt_1_21, // sfix19_En18 
    input [18:0] Wgt_1_22, // sfix19_En18 
    input [18:0] Wgt_1_23, // sfix19_En18 
    input [18:0] Wgt_1_24, // sfix19_En18 
    input [18:0] Wgt_1_25, // sfix19_En18 
    input [18:0] Wgt_1_26, // sfix19_En18 
    input [18:0] Wgt_1_27, // sfix19_En18 
    input [18:0] Wgt_1_28, // sfix19_En18 
    input [18:0] Wgt_1_29, // sfix19_En18 
    input [18:0] Wgt_1_30, // sfix19_En18 
    input [18:0] Wgt_1_31, // sfix19_En18 
    input [18:0] Wgt_1_32, // sfix19_En18 
    input [18:0] Wgt_1_33, // sfix19_En18 
    input [18:0] Wgt_1_34, // sfix19_En18 
    input [18:0] Wgt_1_35, // sfix19_En18 
    input [18:0] Wgt_1_36, // sfix19_En18 
    input [18:0] Wgt_1_37, // sfix19_En18 
    input [18:0] Wgt_1_38, // sfix19_En18 
    input [18:0] Wgt_1_39, // sfix19_En18 
    input [18:0] Wgt_1_40, // sfix19_En18 
    input [18:0] Wgt_1_41, // sfix19_En18 
    input [18:0] Wgt_1_42, // sfix19_En18 
    input [18:0] Wgt_1_43, // sfix19_En18 
    input [18:0] Wgt_1_44, // sfix19_En18 
    input [18:0] Wgt_1_45, // sfix19_En18 
    input [18:0] Wgt_1_46, // sfix19_En18 
    input [18:0] Wgt_1_47, // sfix19_En18 
    input [18:0] Wgt_1_48, // sfix19_En18 
    input [18:0] Wgt_1_49, // sfix19_En18 
    input [18:0] Wgt_1_50, // sfix19_En18 
    input [18:0] Wgt_1_51, // sfix19_En18 
    input [18:0] Wgt_1_52, // sfix19_En18 
    input [18:0] Wgt_1_53, // sfix19_En18 
    input [18:0] Wgt_1_54, // sfix19_En18 
    input [18:0] Wgt_1_55, // sfix19_En18 
    input [18:0] Wgt_1_56, // sfix19_En18 
    input [18:0] Wgt_1_57, // sfix19_En18 
    input [18:0] Wgt_1_58, // sfix19_En18 
    input [18:0] Wgt_1_59, // sfix19_En18 
    input [18:0] Wgt_1_60, // sfix19_En18 
    input [18:0] Wgt_1_61, // sfix19_En18 
    input [18:0] Wgt_1_62, // sfix19_En18 
    input [18:0] Wgt_1_63, // sfix19_En18 
    input [18:0] Wgt_1_64, // sfix19_En18 
    input [18:0] Wgt_1_65, // sfix19_En18 
    input [18:0] Wgt_1_66, // sfix19_En18 
    input [18:0] Wgt_1_67, // sfix19_En18 
    input [18:0] Wgt_1_68, // sfix19_En18 
    input [18:0] Wgt_1_69, // sfix19_En18 
    input [18:0] Wgt_1_70, // sfix19_En18 
    input [18:0] Wgt_1_71, // sfix19_En18 
    input [18:0] Wgt_1_72, // sfix19_En18 
    input [18:0] Wgt_1_73, // sfix19_En18 
    input [18:0] Wgt_1_74, // sfix19_En18 
    input [18:0] Wgt_1_75, // sfix19_En18 
    input [18:0] Wgt_1_76, // sfix19_En18 
    input [18:0] Wgt_1_77, // sfix19_En18 
    input [18:0] Wgt_1_78, // sfix19_En18 
    input [18:0] Wgt_1_79, // sfix19_En18 
    input [18:0] Wgt_1_80, // sfix19_En18 
    input [18:0] Wgt_1_81, // sfix19_En18 
    input [18:0] Wgt_1_82, // sfix19_En18 
    input [18:0] Wgt_1_83, // sfix19_En18 
    input [18:0] Wgt_1_84, // sfix19_En18 
    input [18:0] Wgt_1_85, // sfix19_En18 
    input [18:0] Wgt_1_86, // sfix19_En18 
    input [18:0] Wgt_1_87, // sfix19_En18 
    input [18:0] Wgt_1_88, // sfix19_En18 
    input [18:0] Wgt_1_89, // sfix19_En18 
    input [18:0] Wgt_1_90, // sfix19_En18 
    input [18:0] Wgt_1_91, // sfix19_En18 
    input [18:0] Wgt_1_92, // sfix19_En18 
    input [18:0] Wgt_1_93, // sfix19_En18 
    input [18:0] Wgt_1_94, // sfix19_En18 
    input [18:0] Wgt_1_95, // sfix19_En18 
    input [18:0] Wgt_1_96, // sfix19_En18 
    input [18:0] Wgt_1_97, // sfix19_En18 
    input [18:0] Wgt_1_98, // sfix19_En18 
    input [18:0] Wgt_1_99, // sfix19_En18 
    input [18:0] Wgt_1_100, // sfix19_En18 
    input [18:0] Wgt_1_101, // sfix19_En18 
    input [18:0] Wgt_1_102, // sfix19_En18 
    input [18:0] Wgt_1_103, // sfix19_En18 
    input [18:0] Wgt_1_104, // sfix19_En18 
    input [18:0] Wgt_1_105, // sfix19_En18 
    input [18:0] Wgt_1_106, // sfix19_En18 
    input [18:0] Wgt_1_107, // sfix19_En18 
    input [18:0] Wgt_1_108, // sfix19_En18 
    input [18:0] Wgt_1_109, // sfix19_En18 
    input [18:0] Wgt_1_110, // sfix19_En18 
    input [18:0] Wgt_1_111, // sfix19_En18 
    input [18:0] Wgt_1_112, // sfix19_En18 
    input [18:0] Wgt_1_113, // sfix19_En18 
    input [18:0] Wgt_1_114, // sfix19_En18 
    input [18:0] Wgt_1_115, // sfix19_En18 
    input [18:0] Wgt_1_116, // sfix19_En18 
    input [18:0] Wgt_1_117, // sfix19_En18 
    input [18:0] Wgt_1_118, // sfix19_En18 
    input [18:0] Wgt_1_119, // sfix19_En18 
    input [18:0] Wgt_1_120, // sfix19_En18 
    input [18:0] Wgt_1_121, // sfix19_En18 
    input [18:0] Wgt_1_122, // sfix19_En18 
    input [18:0] Wgt_1_123, // sfix19_En18 
    input [18:0] Wgt_1_124, // sfix19_En18 
    input [18:0] Wgt_1_125, // sfix19_En18 
    input [18:0] Wgt_1_126, // sfix19_En18 
    input [18:0] Wgt_1_127, // sfix19_En18 
    input [18:0] Wgt_1_128, // sfix19_En18 
    input [18:0] Wgt_1_129, // sfix19_En18 
    input [18:0] Wgt_1_130, // sfix19_En18 
    input [18:0] Wgt_1_131, // sfix19_En18 
    input [18:0] Wgt_1_132, // sfix19_En18 
    input [18:0] Wgt_1_133, // sfix19_En18 
    input [18:0] Wgt_1_134, // sfix19_En18 
    input [18:0] Wgt_1_135, // sfix19_En18 
    input [18:0] Wgt_1_136, // sfix19_En18 
    input [18:0] Wgt_1_137, // sfix19_En18 
    input [18:0] Wgt_1_138, // sfix19_En18 
    input [18:0] Wgt_1_139, // sfix19_En18 
    input [18:0] Wgt_1_140, // sfix19_En18 
    input [18:0] Wgt_1_141, // sfix19_En18 
    input [18:0] Wgt_1_142, // sfix19_En18 
    input [18:0] Wgt_1_143, // sfix19_En18 
    input [18:0] Wgt_1_144, // sfix19_En18 
    input [18:0] Wgt_1_145, // sfix19_En18 
    input [18:0] Wgt_1_146, // sfix19_En18 
    input [18:0] Wgt_1_147, // sfix19_En18 
    input [18:0] Wgt_1_148, // sfix19_En18 
    input [18:0] Wgt_1_149, // sfix19_En18 
    input [18:0] Wgt_1_150, // sfix19_En18 
    input [18:0] Wgt_1_151, // sfix19_En18 
    input [18:0] Wgt_1_152, // sfix19_En18 
    input [18:0] Wgt_1_153, // sfix19_En18 
    input [18:0] Wgt_1_154, // sfix19_En18 
    input [18:0] Wgt_1_155, // sfix19_En18 
    input [18:0] Wgt_1_156, // sfix19_En18 
    input [18:0] Wgt_1_157, // sfix19_En18 
    input [18:0] Wgt_1_158, // sfix19_En18 
    input [18:0] Wgt_1_159, // sfix19_En18 
    input [18:0] Wgt_1_160, // sfix19_En18 
    input [18:0] Wgt_1_161, // sfix19_En18 
    input [18:0] Wgt_1_162, // sfix19_En18 
    input [18:0] Wgt_1_163, // sfix19_En18 
    input [18:0] Wgt_1_164, // sfix19_En18 
    input [18:0] Wgt_1_165, // sfix19_En18 
    input [18:0] Wgt_1_166, // sfix19_En18 
    input [18:0] Wgt_1_167, // sfix19_En18 
    input [18:0] Wgt_1_168, // sfix19_En18 
    input [18:0] Wgt_1_169, // sfix19_En18 
    input [18:0] Wgt_1_170, // sfix19_En18 
    input [18:0] Wgt_1_171, // sfix19_En18 
    input [18:0] Wgt_1_172, // sfix19_En18 
    input [18:0] Wgt_1_173, // sfix19_En18 
    input [18:0] Wgt_1_174, // sfix19_En18 
    input [18:0] Wgt_1_175, // sfix19_En18 
    input [18:0] Wgt_1_176, // sfix19_En18 
    input [18:0] Wgt_1_177, // sfix19_En18 
    input [18:0] Wgt_1_178, // sfix19_En18 
    input [18:0] Wgt_1_179, // sfix19_En18 
    input [18:0] Wgt_1_180, // sfix19_En18 
    input [18:0] Wgt_1_181, // sfix19_En18 
    input [18:0] Wgt_1_182, // sfix19_En18 
    input [18:0] Wgt_1_183, // sfix19_En18 
    input [18:0] Wgt_1_184, // sfix19_En18 
    input [18:0] Wgt_1_185, // sfix19_En18 
    input [18:0] Wgt_1_186, // sfix19_En18 
    input [18:0] Wgt_1_187, // sfix19_En18 
    input [18:0] Wgt_1_188, // sfix19_En18 
    input [18:0] Wgt_1_189, // sfix19_En18 
    input [18:0] Wgt_1_190, // sfix19_En18 
    input [18:0] Wgt_1_191, // sfix19_En18 
    input [18:0] Wgt_1_192, // sfix19_En18 
    input [18:0] Wgt_1_193, // sfix19_En18 
    input [18:0] Wgt_1_194, // sfix19_En18 
    input [18:0] Wgt_1_195, // sfix19_En18 
    input [18:0] Wgt_1_196, // sfix19_En18 
    input [18:0] Wgt_1_197, // sfix19_En18 
    input [18:0] Wgt_1_198, // sfix19_En18 
    input [18:0] Wgt_1_199, // sfix19_En18 
    input [18:0] Wgt_1_200, // sfix19_En18 
    input [18:0] Wgt_1_201, // sfix19_En18 
    input [18:0] Wgt_1_202, // sfix19_En18 
    input [18:0] Wgt_1_203, // sfix19_En18 
    input [18:0] Wgt_1_204, // sfix19_En18 
    input [18:0] Wgt_1_205, // sfix19_En18 
    input [18:0] Wgt_1_206, // sfix19_En18 
    input [18:0] Wgt_1_207, // sfix19_En18 
    input [18:0] Wgt_1_208, // sfix19_En18 
    input [18:0] Wgt_1_209, // sfix19_En18 
    input [18:0] Wgt_1_210, // sfix19_En18 
    input [18:0] Wgt_1_211, // sfix19_En18 
    input [18:0] Wgt_1_212, // sfix19_En18 
    input [18:0] Wgt_1_213, // sfix19_En18 
    input [18:0] Wgt_1_214, // sfix19_En18 
    input [18:0] Wgt_1_215, // sfix19_En18 
    input [18:0] Wgt_1_216, // sfix19_En18 
    input [18:0] Wgt_1_217, // sfix19_En18 
    input [18:0] Wgt_1_218, // sfix19_En18 
    input [18:0] Wgt_1_219, // sfix19_En18 
    input [18:0] Wgt_1_220, // sfix19_En18 
    input [18:0] Wgt_1_221, // sfix19_En18 
    input [18:0] Wgt_1_222, // sfix19_En18 
    input [18:0] Wgt_1_223, // sfix19_En18 
    input [18:0] Wgt_1_224, // sfix19_En18 
    input [18:0] Wgt_1_225, // sfix19_En18 
    input [18:0] Wgt_1_226, // sfix19_En18 
    input [18:0] Wgt_1_227, // sfix19_En18 
    input [18:0] Wgt_1_228, // sfix19_En18 
    input [18:0] Wgt_1_229, // sfix19_En18 
    input [18:0] Wgt_1_230, // sfix19_En18 
    input [18:0] Wgt_1_231, // sfix19_En18 
    input [18:0] Wgt_1_232, // sfix19_En18 
    input [18:0] Wgt_1_233, // sfix19_En18 
    input [18:0] Wgt_1_234, // sfix19_En18 
    input [18:0] Wgt_1_235, // sfix19_En18 
    input [18:0] Wgt_1_236, // sfix19_En18 
    input [18:0] Wgt_1_237, // sfix19_En18 
    input [18:0] Wgt_1_238, // sfix19_En18 
    input [18:0] Wgt_1_239, // sfix19_En18 
    input [18:0] Wgt_1_240, // sfix19_En18 
    input [18:0] Wgt_1_241, // sfix19_En18 
    input [18:0] Wgt_1_242, // sfix19_En18 
    input [18:0] Wgt_1_243, // sfix19_En18 
    input [18:0] Wgt_1_244, // sfix19_En18 
    input [18:0] Wgt_1_245, // sfix19_En18 
    input [18:0] Wgt_1_246, // sfix19_En18 
    input [18:0] Wgt_1_247, // sfix19_En18 
    input [18:0] Wgt_1_248, // sfix19_En18 
    input [18:0] Wgt_1_249, // sfix19_En18 
    input [18:0] Wgt_1_250, // sfix19_En18 
    input [18:0] Wgt_1_251, // sfix19_En18 
    input [18:0] Wgt_1_252, // sfix19_En18 
    input [18:0] Wgt_1_253, // sfix19_En18 
    input [18:0] Wgt_1_254, // sfix19_En18 
    input [18:0] Wgt_1_255, // sfix19_En18 
    input [18:0] Wgt_1_256, // sfix19_En18 
    input [18:0] Wgt_1_257, // sfix19_En18 
    input [18:0] Wgt_1_258, // sfix19_En18 
    input [18:0] Wgt_1_259, // sfix19_En18 
    input [18:0] Wgt_1_260, // sfix19_En18 
    input [18:0] Wgt_1_261, // sfix19_En18 
    input [18:0] Wgt_1_262, // sfix19_En18 
    input [18:0] Wgt_1_263, // sfix19_En18 
    input [18:0] Wgt_1_264, // sfix19_En18 
    input [18:0] Wgt_1_265, // sfix19_En18 
    input [18:0] Wgt_1_266, // sfix19_En18 
    input [18:0] Wgt_1_267, // sfix19_En18 
    input [18:0] Wgt_1_268, // sfix19_En18 
    input [18:0] Wgt_1_269, // sfix19_En18 
    input [18:0] Wgt_1_270, // sfix19_En18 
    input [18:0] Wgt_1_271, // sfix19_En18 
    input [18:0] Wgt_1_272, // sfix19_En18 
    input [18:0] Wgt_1_273, // sfix19_En18 
    input [18:0] Wgt_1_274, // sfix19_En18 
    input [18:0] Wgt_1_275, // sfix19_En18 
    input [18:0] Wgt_1_276, // sfix19_En18 
    input [18:0] Wgt_1_277, // sfix19_En18 
    input [18:0] Wgt_1_278, // sfix19_En18 
    input [18:0] Wgt_1_279, // sfix19_En18 
    input [18:0] Wgt_1_280, // sfix19_En18 
    input [18:0] Wgt_1_281, // sfix19_En18 
    input [18:0] Wgt_1_282, // sfix19_En18 
    input [18:0] Wgt_1_283, // sfix19_En18 
    input [18:0] Wgt_1_284, // sfix19_En18 
    input [18:0] Wgt_1_285, // sfix19_En18 
    input [18:0] Wgt_1_286, // sfix19_En18 
    input [18:0] Wgt_1_287, // sfix19_En18 
    input [18:0] Wgt_1_288, // sfix19_En18 
    input [18:0] Wgt_1_289, // sfix19_En18 
    input [18:0] Wgt_1_290, // sfix19_En18 
    input [18:0] Wgt_1_291, // sfix19_En18 
    input [18:0] Wgt_1_292, // sfix19_En18 
    input [18:0] Wgt_1_293, // sfix19_En18 
    input [18:0] Wgt_1_294, // sfix19_En18 
    input [18:0] Wgt_1_295, // sfix19_En18 
    input [18:0] Wgt_1_296, // sfix19_En18 
    input [18:0] Wgt_1_297, // sfix19_En18 
    input [18:0] Wgt_1_298, // sfix19_En18 
    input [18:0] Wgt_1_299, // sfix19_En18 
    input [18:0] Wgt_1_300, // sfix19_En18 
    input [18:0] Wgt_1_301, // sfix19_En18 
    input [18:0] Wgt_1_302, // sfix19_En18 
    input [18:0] Wgt_1_303, // sfix19_En18 
    input [18:0] Wgt_1_304, // sfix19_En18 
    input [18:0] Wgt_1_305, // sfix19_En18 
    input [18:0] Wgt_1_306, // sfix19_En18 
    input [18:0] Wgt_1_307, // sfix19_En18 
    input [18:0] Wgt_1_308, // sfix19_En18 
    input [18:0] Wgt_1_309, // sfix19_En18 
    input [18:0] Wgt_1_310, // sfix19_En18 
    input [18:0] Wgt_1_311, // sfix19_En18 
    input [18:0] Wgt_1_312, // sfix19_En18 
    input [18:0] Wgt_1_313, // sfix19_En18 
    input [18:0] Wgt_1_314, // sfix19_En18 
    input [18:0] Wgt_1_315, // sfix19_En18 
    input [18:0] Wgt_1_316, // sfix19_En18 
    input [18:0] Wgt_1_317, // sfix19_En18 
    input [18:0] Wgt_1_318, // sfix19_En18 
    input [18:0] Wgt_1_319, // sfix19_En18 
    input [18:0] Wgt_1_320, // sfix19_En18 
    input [18:0] Wgt_1_321, // sfix19_En18 
    input [18:0] Wgt_1_322, // sfix19_En18 
    input [18:0] Wgt_1_323, // sfix19_En18 
    input [18:0] Wgt_1_324, // sfix19_En18 
    input [18:0] Wgt_1_325, // sfix19_En18 
    input [18:0] Wgt_1_326, // sfix19_En18 
    input [18:0] Wgt_1_327, // sfix19_En18 
    input [18:0] Wgt_1_328, // sfix19_En18 
    input [18:0] Wgt_1_329, // sfix19_En18 
    input [18:0] Wgt_1_330, // sfix19_En18 
    input [18:0] Wgt_1_331, // sfix19_En18 
    input [18:0] Wgt_1_332, // sfix19_En18 
    input [18:0] Wgt_1_333, // sfix19_En18 
    input [18:0] Wgt_1_334, // sfix19_En18 
    input [18:0] Wgt_1_335, // sfix19_En18 
    input [18:0] Wgt_1_336, // sfix19_En18 
    input [18:0] Wgt_1_337, // sfix19_En18 
    input [18:0] Wgt_1_338, // sfix19_En18 
    input [18:0] Wgt_1_339, // sfix19_En18 
    input [18:0] Wgt_1_340, // sfix19_En18 
    input [18:0] Wgt_1_341, // sfix19_En18 
    input [18:0] Wgt_1_342, // sfix19_En18 
    input [18:0] Wgt_1_343, // sfix19_En18 
    input [18:0] Wgt_1_344, // sfix19_En18 
    input [18:0] Wgt_1_345, // sfix19_En18 
    input [18:0] Wgt_1_346, // sfix19_En18 
    input [18:0] Wgt_1_347, // sfix19_En18 
    input [18:0] Wgt_1_348, // sfix19_En18 
    input [18:0] Wgt_1_349, // sfix19_En18 
    input [18:0] Wgt_1_350, // sfix19_En18 
    input [18:0] Wgt_1_351, // sfix19_En18 
    input [18:0] Wgt_1_352, // sfix19_En18 
    input [18:0] Wgt_1_353, // sfix19_En18 
    input [18:0] Wgt_1_354, // sfix19_En18 
    input [18:0] Wgt_1_355, // sfix19_En18 
    input [18:0] Wgt_1_356, // sfix19_En18 
    input [18:0] Wgt_1_357, // sfix19_En18 
    input [18:0] Wgt_1_358, // sfix19_En18 
    input [18:0] Wgt_1_359, // sfix19_En18 
    input [18:0] Wgt_1_360, // sfix19_En18 
    input [18:0] Wgt_1_361, // sfix19_En18 
    input [18:0] Wgt_1_362, // sfix19_En18 
    input [18:0] Wgt_1_363, // sfix19_En18 
    input [18:0] Wgt_1_364, // sfix19_En18 
    input [18:0] Wgt_1_365, // sfix19_En18 
    input [18:0] Wgt_1_366, // sfix19_En18 
    input [18:0] Wgt_1_367, // sfix19_En18 
    input [18:0] Wgt_1_368, // sfix19_En18 
    input [18:0] Wgt_1_369, // sfix19_En18 
    input [18:0] Wgt_1_370, // sfix19_En18 
    input [18:0] Wgt_1_371, // sfix19_En18 
    input [18:0] Wgt_1_372, // sfix19_En18 
    input [18:0] Wgt_1_373, // sfix19_En18 
    input [18:0] Wgt_1_374, // sfix19_En18 
    input [18:0] Wgt_1_375, // sfix19_En18 
    input [18:0] Wgt_1_376, // sfix19_En18 
    input [18:0] Wgt_1_377, // sfix19_En18 
    input [18:0] Wgt_1_378, // sfix19_En18 
    input [18:0] Wgt_1_379, // sfix19_En18 
    input [18:0] Wgt_1_380, // sfix19_En18 
    input [18:0] Wgt_1_381, // sfix19_En18 
    input [18:0] Wgt_1_382, // sfix19_En18 
    input [18:0] Wgt_1_383, // sfix19_En18 
    input [18:0] Wgt_1_384, // sfix19_En18 
    input [18:0] Wgt_1_385, // sfix19_En18 
    input [18:0] Wgt_1_386, // sfix19_En18 
    input [18:0] Wgt_1_387, // sfix19_En18 
    input [18:0] Wgt_1_388, // sfix19_En18 
    input [18:0] Wgt_1_389, // sfix19_En18 
    input [18:0] Wgt_1_390, // sfix19_En18 
    input [18:0] Wgt_1_391, // sfix19_En18 
    input [18:0] Wgt_1_392, // sfix19_En18 
    input [18:0] Wgt_1_393, // sfix19_En18 
    input [18:0] Wgt_1_394, // sfix19_En18 
    input [18:0] Wgt_1_395, // sfix19_En18 
    input [18:0] Wgt_1_396, // sfix19_En18 
    input [18:0] Wgt_1_397, // sfix19_En18 
    input [18:0] Wgt_1_398, // sfix19_En18 
    input [18:0] Wgt_1_399, // sfix19_En18 
    input [18:0] Wgt_1_400, // sfix19_En18 
    input [18:0] Wgt_1_401, // sfix19_En18 
    input [18:0] Wgt_1_402, // sfix19_En18 
    input [18:0] Wgt_1_403, // sfix19_En18 
    input [18:0] Wgt_1_404, // sfix19_En18 
    input [18:0] Wgt_1_405, // sfix19_En18 
    input [18:0] Wgt_1_406, // sfix19_En18 
    input [18:0] Wgt_1_407, // sfix19_En18 
    input [18:0] Wgt_1_408, // sfix19_En18 
    input [18:0] Wgt_1_409, // sfix19_En18 
    input [18:0] Wgt_1_410, // sfix19_En18 
    input [18:0] Wgt_1_411, // sfix19_En18 
    input [18:0] Wgt_1_412, // sfix19_En18 
    input [18:0] Wgt_1_413, // sfix19_En18 
    input [18:0] Wgt_1_414, // sfix19_En18 
    input [18:0] Wgt_1_415, // sfix19_En18 
    input [18:0] Wgt_1_416, // sfix19_En18 
    input [18:0] Wgt_1_417, // sfix19_En18 
    input [18:0] Wgt_1_418, // sfix19_En18 
    input [18:0] Wgt_1_419, // sfix19_En18 
    input [18:0] Wgt_1_420, // sfix19_En18 
    input [18:0] Wgt_1_421, // sfix19_En18 
    input [18:0] Wgt_1_422, // sfix19_En18 
    input [18:0] Wgt_1_423, // sfix19_En18 
    input [18:0] Wgt_1_424, // sfix19_En18 
    input [18:0] Wgt_1_425, // sfix19_En18 
    input [18:0] Wgt_1_426, // sfix19_En18 
    input [18:0] Wgt_1_427, // sfix19_En18 
    input [18:0] Wgt_1_428, // sfix19_En18 
    input [18:0] Wgt_1_429, // sfix19_En18 
    input [18:0] Wgt_1_430, // sfix19_En18 
    input [18:0] Wgt_1_431, // sfix19_En18 
    input [18:0] Wgt_1_432, // sfix19_En18 
    input [18:0] Wgt_1_433, // sfix19_En18 
    input [18:0] Wgt_1_434, // sfix19_En18 
    input [18:0] Wgt_1_435, // sfix19_En18 
    input [18:0] Wgt_1_436, // sfix19_En18 
    input [18:0] Wgt_1_437, // sfix19_En18 
    input [18:0] Wgt_1_438, // sfix19_En18 
    input [18:0] Wgt_1_439, // sfix19_En18 
    input [18:0] Wgt_1_440, // sfix19_En18 
    input [18:0] Wgt_1_441, // sfix19_En18 
    input [18:0] Wgt_1_442, // sfix19_En18 
    input [18:0] Wgt_1_443, // sfix19_En18 
    input [18:0] Wgt_1_444, // sfix19_En18 
    input [18:0] Wgt_1_445, // sfix19_En18 
    input [18:0] Wgt_1_446, // sfix19_En18 
    input [18:0] Wgt_1_447, // sfix19_En18 
    input [18:0] Wgt_1_448, // sfix19_En18 
    input [18:0] Wgt_1_449, // sfix19_En18 
    input [18:0] Wgt_1_450, // sfix19_En18 
    input [18:0] Wgt_1_451, // sfix19_En18 
    input [18:0] Wgt_1_452, // sfix19_En18 
    input [18:0] Wgt_1_453, // sfix19_En18 
    input [18:0] Wgt_1_454, // sfix19_En18 
    input [18:0] Wgt_1_455, // sfix19_En18 
    input [18:0] Wgt_1_456, // sfix19_En18 
    input [18:0] Wgt_1_457, // sfix19_En18 
    input [18:0] Wgt_1_458, // sfix19_En18 
    input [18:0] Wgt_1_459, // sfix19_En18 
    input [18:0] Wgt_1_460, // sfix19_En18 
    input [18:0] Wgt_1_461, // sfix19_En18 
    input [18:0] Wgt_1_462, // sfix19_En18 
    input [18:0] Wgt_1_463, // sfix19_En18 
    input [18:0] Wgt_1_464, // sfix19_En18 
    input [18:0] Wgt_1_465, // sfix19_En18 
    input [18:0] Wgt_1_466, // sfix19_En18 
    input [18:0] Wgt_1_467, // sfix19_En18 
    input [18:0] Wgt_1_468, // sfix19_En18 
    input [18:0] Wgt_1_469, // sfix19_En18 
    input [18:0] Wgt_1_470, // sfix19_En18 
    input [18:0] Wgt_1_471, // sfix19_En18 
    input [18:0] Wgt_1_472, // sfix19_En18 
    input [18:0] Wgt_1_473, // sfix19_En18 
    input [18:0] Wgt_1_474, // sfix19_En18 
    input [18:0] Wgt_1_475, // sfix19_En18 
    input [18:0] Wgt_1_476, // sfix19_En18 
    input [18:0] Wgt_1_477, // sfix19_En18 
    input [18:0] Wgt_1_478, // sfix19_En18 
    input [18:0] Wgt_1_479, // sfix19_En18 
    input [18:0] Wgt_1_480, // sfix19_En18 
    input [18:0] Wgt_1_481, // sfix19_En18 
    input [18:0] Wgt_1_482, // sfix19_En18 
    input [18:0] Wgt_1_483, // sfix19_En18 
    input [18:0] Wgt_1_484, // sfix19_En18 
    input [18:0] Wgt_1_485, // sfix19_En18 
    input [18:0] Wgt_1_486, // sfix19_En18 
    input [18:0] Wgt_1_487, // sfix19_En18 
    input [18:0] Wgt_1_488, // sfix19_En18 
    input [18:0] Wgt_1_489, // sfix19_En18 
    input [18:0] Wgt_1_490, // sfix19_En18 
    input [18:0] Wgt_1_491, // sfix19_En18 
    input [18:0] Wgt_1_492, // sfix19_En18 
    input [18:0] Wgt_1_493, // sfix19_En18 
    input [18:0] Wgt_1_494, // sfix19_En18 
    input [18:0] Wgt_1_495, // sfix19_En18 
    input [18:0] Wgt_1_496, // sfix19_En18 
    input [18:0] Wgt_1_497, // sfix19_En18 
    input [18:0] Wgt_1_498, // sfix19_En18 
    input [18:0] Wgt_1_499, // sfix19_En18 
    input [18:0] Wgt_1_500, // sfix19_En18 
    input [18:0] Wgt_1_501, // sfix19_En18 
    input [18:0] Wgt_1_502, // sfix19_En18 
    input [18:0] Wgt_1_503, // sfix19_En18 
    input [18:0] Wgt_1_504, // sfix19_En18 
    input [18:0] Wgt_1_505, // sfix19_En18 
    input [18:0] Wgt_1_506, // sfix19_En18 
    input [18:0] Wgt_1_507, // sfix19_En18 
    input [18:0] Wgt_1_508, // sfix19_En18 
    input [18:0] Wgt_1_509, // sfix19_En18 
    input [18:0] Wgt_1_510, // sfix19_En18 
    input [18:0] Wgt_1_511, // sfix19_En18 
    input [18:0] Wgt_1_512, // sfix19_En18 
    input [18:0] Wgt_1_513, // sfix19_En18 
    input [18:0] Wgt_1_514, // sfix19_En18 
    input [18:0] Wgt_1_515, // sfix19_En18 
    input [18:0] Wgt_1_516, // sfix19_En18 
    input [18:0] Wgt_1_517, // sfix19_En18 
    input [18:0] Wgt_1_518, // sfix19_En18 
    input [18:0] Wgt_1_519, // sfix19_En18 
    input [18:0] Wgt_1_520, // sfix19_En18 
    input [18:0] Wgt_1_521, // sfix19_En18 
    input [18:0] Wgt_1_522, // sfix19_En18 
    input [18:0] Wgt_1_523, // sfix19_En18 
    input [18:0] Wgt_1_524, // sfix19_En18 
    input [18:0] Wgt_1_525, // sfix19_En18 
    input [18:0] Wgt_1_526, // sfix19_En18 
    input [18:0] Wgt_1_527, // sfix19_En18 
    input [18:0] Wgt_1_528, // sfix19_En18 
    input [18:0] Wgt_1_529, // sfix19_En18 
    input [18:0] Wgt_1_530, // sfix19_En18 
    input [18:0] Wgt_1_531, // sfix19_En18 
    input [18:0] Wgt_1_532, // sfix19_En18 
    input [18:0] Wgt_1_533, // sfix19_En18 
    input [18:0] Wgt_1_534, // sfix19_En18 
    input [18:0] Wgt_1_535, // sfix19_En18 
    input [18:0] Wgt_1_536, // sfix19_En18 
    input [18:0] Wgt_1_537, // sfix19_En18 
    input [18:0] Wgt_1_538, // sfix19_En18 
    input [18:0] Wgt_1_539, // sfix19_En18 
    input [18:0] Wgt_1_540, // sfix19_En18 
    input [18:0] Wgt_1_541, // sfix19_En18 
    input [18:0] Wgt_1_542, // sfix19_En18 
    input [18:0] Wgt_1_543, // sfix19_En18 
    input [18:0] Wgt_1_544, // sfix19_En18 
    input [18:0] Wgt_1_545, // sfix19_En18 
    input [18:0] Wgt_1_546, // sfix19_En18 
    input [18:0] Wgt_1_547, // sfix19_En18 
    input [18:0] Wgt_1_548, // sfix19_En18 
    input [18:0] Wgt_1_549, // sfix19_En18 
    input [18:0] Wgt_1_550, // sfix19_En18 
    input [18:0] Wgt_1_551, // sfix19_En18 
    input [18:0] Wgt_1_552, // sfix19_En18 
    input [18:0] Wgt_1_553, // sfix19_En18 
    input [18:0] Wgt_1_554, // sfix19_En18 
    input [18:0] Wgt_1_555, // sfix19_En18 
    input [18:0] Wgt_1_556, // sfix19_En18 
    input [18:0] Wgt_1_557, // sfix19_En18 
    input [18:0] Wgt_1_558, // sfix19_En18 
    input [18:0] Wgt_1_559, // sfix19_En18 
    input [18:0] Wgt_1_560, // sfix19_En18 
    input [18:0] Wgt_1_561, // sfix19_En18 
    input [18:0] Wgt_1_562, // sfix19_En18 
    input [18:0] Wgt_1_563, // sfix19_En18 
    input [18:0] Wgt_1_564, // sfix19_En18 
    input [18:0] Wgt_1_565, // sfix19_En18 
    input [18:0] Wgt_1_566, // sfix19_En18 
    input [18:0] Wgt_1_567, // sfix19_En18 
    input [18:0] Wgt_1_568, // sfix19_En18 
    input [18:0] Wgt_1_569, // sfix19_En18 
    input [18:0] Wgt_1_570, // sfix19_En18 
    input [18:0] Wgt_1_571, // sfix19_En18 
    input [18:0] Wgt_1_572, // sfix19_En18 
    input [18:0] Wgt_1_573, // sfix19_En18 
    input [18:0] Wgt_1_574, // sfix19_En18 
    input [18:0] Wgt_1_575, // sfix19_En18 
    input [18:0] Wgt_1_576, // sfix19_En18 
    input [18:0] Wgt_1_577, // sfix19_En18 
    input [18:0] Wgt_1_578, // sfix19_En18 
    input [18:0] Wgt_1_579, // sfix19_En18 
    input [18:0] Wgt_1_580, // sfix19_En18 
    input [18:0] Wgt_1_581, // sfix19_En18 
    input [18:0] Wgt_1_582, // sfix19_En18 
    input [18:0] Wgt_1_583, // sfix19_En18 
    input [18:0] Wgt_1_584, // sfix19_En18 
    input [18:0] Wgt_1_585, // sfix19_En18 
    input [18:0] Wgt_1_586, // sfix19_En18 
    input [18:0] Wgt_1_587, // sfix19_En18 
    input [18:0] Wgt_1_588, // sfix19_En18 
    input [18:0] Wgt_1_589, // sfix19_En18 
    input [18:0] Wgt_1_590, // sfix19_En18 
    input [18:0] Wgt_1_591, // sfix19_En18 
    input [18:0] Wgt_1_592, // sfix19_En18 
    input [18:0] Wgt_1_593, // sfix19_En18 
    input [18:0] Wgt_1_594, // sfix19_En18 
    input [18:0] Wgt_1_595, // sfix19_En18 
    input [18:0] Wgt_1_596, // sfix19_En18 
    input [18:0] Wgt_1_597, // sfix19_En18 
    input [18:0] Wgt_1_598, // sfix19_En18 
    input [18:0] Wgt_1_599, // sfix19_En18 
    input [18:0] Wgt_1_600, // sfix19_En18 
    input [18:0] Wgt_1_601, // sfix19_En18 
    input [18:0] Wgt_1_602, // sfix19_En18 
    input [18:0] Wgt_1_603, // sfix19_En18 
    input [18:0] Wgt_1_604, // sfix19_En18 
    input [18:0] Wgt_1_605, // sfix19_En18 
    input [18:0] Wgt_1_606, // sfix19_En18 
    input [18:0] Wgt_1_607, // sfix19_En18 
    input [18:0] Wgt_1_608, // sfix19_En18 
    input [18:0] Wgt_1_609, // sfix19_En18 
    input [18:0] Wgt_1_610, // sfix19_En18 
    input [18:0] Wgt_1_611, // sfix19_En18 
    input [18:0] Wgt_1_612, // sfix19_En18 
    input [18:0] Wgt_1_613, // sfix19_En18 
    input [18:0] Wgt_1_614, // sfix19_En18 
    input [18:0] Wgt_1_615, // sfix19_En18 
    input [18:0] Wgt_1_616, // sfix19_En18 
    input [18:0] Wgt_1_617, // sfix19_En18 
    input [18:0] Wgt_1_618, // sfix19_En18 
    input [18:0] Wgt_1_619, // sfix19_En18 
    input [18:0] Wgt_1_620, // sfix19_En18 
    input [18:0] Wgt_1_621, // sfix19_En18 
    input [18:0] Wgt_1_622, // sfix19_En18 
    input [18:0] Wgt_1_623, // sfix19_En18 
    input [18:0] Wgt_1_624, // sfix19_En18 
    input [18:0] Wgt_1_625, // sfix19_En18 
    input [18:0] Wgt_1_626, // sfix19_En18 
    input [18:0] Wgt_1_627, // sfix19_En18 
    input [18:0] Wgt_1_628, // sfix19_En18 
    input [18:0] Wgt_1_629, // sfix19_En18 
    input [18:0] Wgt_1_630, // sfix19_En18 
    input [18:0] Wgt_1_631, // sfix19_En18 
    input [18:0] Wgt_1_632, // sfix19_En18 
    input [18:0] Wgt_1_633, // sfix19_En18 
    input [18:0] Wgt_1_634, // sfix19_En18 
    input [18:0] Wgt_1_635, // sfix19_En18 
    input [18:0] Wgt_1_636, // sfix19_En18 
    input [18:0] Wgt_1_637, // sfix19_En18 
    input [18:0] Wgt_1_638, // sfix19_En18 
    input [18:0] Wgt_1_639, // sfix19_En18 
    input [18:0] Wgt_1_640, // sfix19_En18 
    input [18:0] Wgt_1_641, // sfix19_En18 
    input [18:0] Wgt_1_642, // sfix19_En18 
    input [18:0] Wgt_1_643, // sfix19_En18 
    input [18:0] Wgt_1_644, // sfix19_En18 
    input [18:0] Wgt_1_645, // sfix19_En18 
    input [18:0] Wgt_1_646, // sfix19_En18 
    input [18:0] Wgt_1_647, // sfix19_En18 
    input [18:0] Wgt_1_648, // sfix19_En18 
    input [18:0] Wgt_1_649, // sfix19_En18 
    input [18:0] Wgt_1_650, // sfix19_En18 
    input [18:0] Wgt_1_651, // sfix19_En18 
    input [18:0] Wgt_1_652, // sfix19_En18 
    input [18:0] Wgt_1_653, // sfix19_En18 
    input [18:0] Wgt_1_654, // sfix19_En18 
    input [18:0] Wgt_1_655, // sfix19_En18 
    input [18:0] Wgt_1_656, // sfix19_En18 
    input [18:0] Wgt_1_657, // sfix19_En18 
    input [18:0] Wgt_1_658, // sfix19_En18 
    input [18:0] Wgt_1_659, // sfix19_En18 
    input [18:0] Wgt_1_660, // sfix19_En18 
    input [18:0] Wgt_1_661, // sfix19_En18 
    input [18:0] Wgt_1_662, // sfix19_En18 
    input [18:0] Wgt_1_663, // sfix19_En18 
    input [18:0] Wgt_1_664, // sfix19_En18 
    input [18:0] Wgt_1_665, // sfix19_En18 
    input [18:0] Wgt_1_666, // sfix19_En18 
    input [18:0] Wgt_1_667, // sfix19_En18 
    input [18:0] Wgt_1_668, // sfix19_En18 
    input [18:0] Wgt_1_669, // sfix19_En18 
    input [18:0] Wgt_1_670, // sfix19_En18 
    input [18:0] Wgt_1_671, // sfix19_En18 
    input [18:0] Wgt_1_672, // sfix19_En18 
    input [18:0] Wgt_1_673, // sfix19_En18 
    input [18:0] Wgt_1_674, // sfix19_En18 
    input [18:0] Wgt_1_675, // sfix19_En18 
    input [18:0] Wgt_1_676, // sfix19_En18 
    input [18:0] Wgt_1_677, // sfix19_En18 
    input [18:0] Wgt_1_678, // sfix19_En18 
    input [18:0] Wgt_1_679, // sfix19_En18 
    input [18:0] Wgt_1_680, // sfix19_En18 
    input [18:0] Wgt_1_681, // sfix19_En18 
    input [18:0] Wgt_1_682, // sfix19_En18 
    input [18:0] Wgt_1_683, // sfix19_En18 
    input [18:0] Wgt_1_684, // sfix19_En18 
    input [18:0] Wgt_1_685, // sfix19_En18 
    input [18:0] Wgt_1_686, // sfix19_En18 
    input [18:0] Wgt_1_687, // sfix19_En18 
    input [18:0] Wgt_1_688, // sfix19_En18 
    input [18:0] Wgt_1_689, // sfix19_En18 
    input [18:0] Wgt_1_690, // sfix19_En18 
    input [18:0] Wgt_1_691, // sfix19_En18 
    input [18:0] Wgt_1_692, // sfix19_En18 
    input [18:0] Wgt_1_693, // sfix19_En18 
    input [18:0] Wgt_1_694, // sfix19_En18 
    input [18:0] Wgt_1_695, // sfix19_En18 
    input [18:0] Wgt_1_696, // sfix19_En18 
    input [18:0] Wgt_1_697, // sfix19_En18 
    input [18:0] Wgt_1_698, // sfix19_En18 
    input [18:0] Wgt_1_699, // sfix19_En18 
    input [18:0] Wgt_1_700, // sfix19_En18 
    input [18:0] Wgt_1_701, // sfix19_En18 
    input [18:0] Wgt_1_702, // sfix19_En18 
    input [18:0] Wgt_1_703, // sfix19_En18 
    input [18:0] Wgt_1_704, // sfix19_En18 
    input [18:0] Wgt_1_705, // sfix19_En18 
    input [18:0] Wgt_1_706, // sfix19_En18 
    input [18:0] Wgt_1_707, // sfix19_En18 
    input [18:0] Wgt_1_708, // sfix19_En18 
    input [18:0] Wgt_1_709, // sfix19_En18 
    input [18:0] Wgt_1_710, // sfix19_En18 
    input [18:0] Wgt_1_711, // sfix19_En18 
    input [18:0] Wgt_1_712, // sfix19_En18 
    input [18:0] Wgt_1_713, // sfix19_En18 
    input [18:0] Wgt_1_714, // sfix19_En18 
    input [18:0] Wgt_1_715, // sfix19_En18 
    input [18:0] Wgt_1_716, // sfix19_En18 
    input [18:0] Wgt_1_717, // sfix19_En18 
    input [18:0] Wgt_1_718, // sfix19_En18 
    input [18:0] Wgt_1_719, // sfix19_En18 
    input [18:0] Wgt_1_720, // sfix19_En18 
    input [18:0] Wgt_1_721, // sfix19_En18 
    input [18:0] Wgt_1_722, // sfix19_En18 
    input [18:0] Wgt_1_723, // sfix19_En18 
    input [18:0] Wgt_1_724, // sfix19_En18 
    input [18:0] Wgt_1_725, // sfix19_En18 
    input [18:0] Wgt_1_726, // sfix19_En18 
    input [18:0] Wgt_1_727, // sfix19_En18 
    input [18:0] Wgt_1_728, // sfix19_En18 
    input [18:0] Wgt_1_729, // sfix19_En18 
    input [18:0] Wgt_1_730, // sfix19_En18 
    input [18:0] Wgt_1_731, // sfix19_En18 
    input [18:0] Wgt_1_732, // sfix19_En18 
    input [18:0] Wgt_1_733, // sfix19_En18 
    input [18:0] Wgt_1_734, // sfix19_En18 
    input [18:0] Wgt_1_735, // sfix19_En18 
    input [18:0] Wgt_1_736, // sfix19_En18 
    input [18:0] Wgt_1_737, // sfix19_En18 
    input [18:0] Wgt_1_738, // sfix19_En18 
    input [18:0] Wgt_1_739, // sfix19_En18 
    input [18:0] Wgt_1_740, // sfix19_En18 
    input [18:0] Wgt_1_741, // sfix19_En18 
    input [18:0] Wgt_1_742, // sfix19_En18 
    input [18:0] Wgt_1_743, // sfix19_En18 
    input [18:0] Wgt_1_744, // sfix19_En18 
    input [18:0] Wgt_1_745, // sfix19_En18 
    input [18:0] Wgt_1_746, // sfix19_En18 
    input [18:0] Wgt_1_747, // sfix19_En18 
    input [18:0] Wgt_1_748, // sfix19_En18 
    input [18:0] Wgt_1_749, // sfix19_En18 
    input [18:0] Wgt_1_750, // sfix19_En18 
    input [18:0] Wgt_1_751, // sfix19_En18 
    input [18:0] Wgt_1_752, // sfix19_En18 
    input [18:0] Wgt_1_753, // sfix19_En18 
    input [18:0] Wgt_1_754, // sfix19_En18 
    input [18:0] Wgt_1_755, // sfix19_En18 
    input [18:0] Wgt_1_756, // sfix19_En18 
    input [18:0] Wgt_1_757, // sfix19_En18 
    input [18:0] Wgt_1_758, // sfix19_En18 
    input [18:0] Wgt_1_759, // sfix19_En18 
    input [18:0] Wgt_1_760, // sfix19_En18 
    input [18:0] Wgt_1_761, // sfix19_En18 
    input [18:0] Wgt_1_762, // sfix19_En18 
    input [18:0] Wgt_1_763, // sfix19_En18 
    input [18:0] Wgt_1_764, // sfix19_En18 
    input [18:0] Wgt_1_765, // sfix19_En18 
    input [18:0] Wgt_1_766, // sfix19_En18 
    input [18:0] Wgt_1_767, // sfix19_En18 
    input [18:0] Wgt_1_768, // sfix19_En18 
    input [18:0] Wgt_1_769, // sfix19_En18 
    input [18:0] Wgt_1_770, // sfix19_En18 
    input [18:0] Wgt_1_771, // sfix19_En18 
    input [18:0] Wgt_1_772, // sfix19_En18 
    input [18:0] Wgt_1_773, // sfix19_En18 
    input [18:0] Wgt_1_774, // sfix19_En18 
    input [18:0] Wgt_1_775, // sfix19_En18 
    input [18:0] Wgt_1_776, // sfix19_En18 
    input [18:0] Wgt_1_777, // sfix19_En18 
    input [18:0] Wgt_1_778, // sfix19_En18 
    input [18:0] Wgt_1_779, // sfix19_En18 
    input [18:0] Wgt_1_780, // sfix19_En18 
    input [18:0] Wgt_1_781, // sfix19_En18 
    input [18:0] Wgt_1_782, // sfix19_En18 
    input [18:0] Wgt_1_783, // sfix19_En18 
    input [18:0] Wgt_1_784, // sfix19_En18 
    input [18:0] Wgt_2_0, // sfix19_En18 
    input [18:0] Wgt_2_1, // sfix19_En18 
    input [18:0] Wgt_2_2, // sfix19_En18 
    input [18:0] Wgt_2_3, // sfix19_En18 
    input [18:0] Wgt_2_4, // sfix19_En18 
    input [18:0] Wgt_2_5, // sfix19_En18 
    input [18:0] Wgt_2_6, // sfix19_En18 
    input [18:0] Wgt_2_7, // sfix19_En18 
    input [18:0] Wgt_2_8, // sfix19_En18 
    input [18:0] Wgt_2_9, // sfix19_En18 
    input [18:0] Wgt_2_10, // sfix19_En18 
    input [18:0] Wgt_2_11, // sfix19_En18 
    input [18:0] Wgt_2_12, // sfix19_En18 
    input [18:0] Wgt_2_13, // sfix19_En18 
    input [18:0] Wgt_2_14, // sfix19_En18 
    input [18:0] Wgt_2_15, // sfix19_En18 
    input [18:0] Wgt_2_16, // sfix19_En18 
    input [18:0] Wgt_2_17, // sfix19_En18 
    input [18:0] Wgt_2_18, // sfix19_En18 
    input [18:0] Wgt_2_19, // sfix19_En18 
    input [18:0] Wgt_2_20, // sfix19_En18 
    input [18:0] Wgt_2_21, // sfix19_En18 
    input [18:0] Wgt_2_22, // sfix19_En18 
    input [18:0] Wgt_2_23, // sfix19_En18 
    input [18:0] Wgt_2_24, // sfix19_En18 
    input [18:0] Wgt_2_25, // sfix19_En18 
    input [18:0] Wgt_2_26, // sfix19_En18 
    input [18:0] Wgt_2_27, // sfix19_En18 
    input [18:0] Wgt_2_28, // sfix19_En18 
    input [18:0] Wgt_2_29, // sfix19_En18 
    input [18:0] Wgt_2_30, // sfix19_En18 
    input [18:0] Wgt_2_31, // sfix19_En18 
    input [18:0] Wgt_2_32, // sfix19_En18 
    input [18:0] Wgt_2_33, // sfix19_En18 
    input [18:0] Wgt_2_34, // sfix19_En18 
    input [18:0] Wgt_2_35, // sfix19_En18 
    input [18:0] Wgt_2_36, // sfix19_En18 
    input [18:0] Wgt_2_37, // sfix19_En18 
    input [18:0] Wgt_2_38, // sfix19_En18 
    input [18:0] Wgt_2_39, // sfix19_En18 
    input [18:0] Wgt_2_40, // sfix19_En18 
    input [18:0] Wgt_2_41, // sfix19_En18 
    input [18:0] Wgt_2_42, // sfix19_En18 
    input [18:0] Wgt_2_43, // sfix19_En18 
    input [18:0] Wgt_2_44, // sfix19_En18 
    input [18:0] Wgt_2_45, // sfix19_En18 
    input [18:0] Wgt_2_46, // sfix19_En18 
    input [18:0] Wgt_2_47, // sfix19_En18 
    input [18:0] Wgt_2_48, // sfix19_En18 
    input [18:0] Wgt_2_49, // sfix19_En18 
    input [18:0] Wgt_2_50, // sfix19_En18 
    input [18:0] Wgt_2_51, // sfix19_En18 
    input [18:0] Wgt_2_52, // sfix19_En18 
    input [18:0] Wgt_2_53, // sfix19_En18 
    input [18:0] Wgt_2_54, // sfix19_En18 
    input [18:0] Wgt_2_55, // sfix19_En18 
    input [18:0] Wgt_2_56, // sfix19_En18 
    input [18:0] Wgt_2_57, // sfix19_En18 
    input [18:0] Wgt_2_58, // sfix19_En18 
    input [18:0] Wgt_2_59, // sfix19_En18 
    input [18:0] Wgt_2_60, // sfix19_En18 
    input [18:0] Wgt_2_61, // sfix19_En18 
    input [18:0] Wgt_2_62, // sfix19_En18 
    input [18:0] Wgt_2_63, // sfix19_En18 
    input [18:0] Wgt_2_64, // sfix19_En18 
    input [18:0] Wgt_2_65, // sfix19_En18 
    input [18:0] Wgt_2_66, // sfix19_En18 
    input [18:0] Wgt_2_67, // sfix19_En18 
    input [18:0] Wgt_2_68, // sfix19_En18 
    input [18:0] Wgt_2_69, // sfix19_En18 
    input [18:0] Wgt_2_70, // sfix19_En18 
    input [18:0] Wgt_2_71, // sfix19_En18 
    input [18:0] Wgt_2_72, // sfix19_En18 
    input [18:0] Wgt_2_73, // sfix19_En18 
    input [18:0] Wgt_2_74, // sfix19_En18 
    input [18:0] Wgt_2_75, // sfix19_En18 
    input [18:0] Wgt_2_76, // sfix19_En18 
    input [18:0] Wgt_2_77, // sfix19_En18 
    input [18:0] Wgt_2_78, // sfix19_En18 
    input [18:0] Wgt_2_79, // sfix19_En18 
    input [18:0] Wgt_2_80, // sfix19_En18 
    input [18:0] Wgt_2_81, // sfix19_En18 
    input [18:0] Wgt_2_82, // sfix19_En18 
    input [18:0] Wgt_2_83, // sfix19_En18 
    input [18:0] Wgt_2_84, // sfix19_En18 
    input [18:0] Wgt_2_85, // sfix19_En18 
    input [18:0] Wgt_2_86, // sfix19_En18 
    input [18:0] Wgt_2_87, // sfix19_En18 
    input [18:0] Wgt_2_88, // sfix19_En18 
    input [18:0] Wgt_2_89, // sfix19_En18 
    input [18:0] Wgt_2_90, // sfix19_En18 
    input [18:0] Wgt_2_91, // sfix19_En18 
    input [18:0] Wgt_2_92, // sfix19_En18 
    input [18:0] Wgt_2_93, // sfix19_En18 
    input [18:0] Wgt_2_94, // sfix19_En18 
    input [18:0] Wgt_2_95, // sfix19_En18 
    input [18:0] Wgt_2_96, // sfix19_En18 
    input [18:0] Wgt_2_97, // sfix19_En18 
    input [18:0] Wgt_2_98, // sfix19_En18 
    input [18:0] Wgt_2_99, // sfix19_En18 
    input [18:0] Wgt_2_100, // sfix19_En18 
    input [18:0] Wgt_2_101, // sfix19_En18 
    input [18:0] Wgt_2_102, // sfix19_En18 
    input [18:0] Wgt_2_103, // sfix19_En18 
    input [18:0] Wgt_2_104, // sfix19_En18 
    input [18:0] Wgt_2_105, // sfix19_En18 
    input [18:0] Wgt_2_106, // sfix19_En18 
    input [18:0] Wgt_2_107, // sfix19_En18 
    input [18:0] Wgt_2_108, // sfix19_En18 
    input [18:0] Wgt_2_109, // sfix19_En18 
    input [18:0] Wgt_2_110, // sfix19_En18 
    input [18:0] Wgt_2_111, // sfix19_En18 
    input [18:0] Wgt_2_112, // sfix19_En18 
    input [18:0] Wgt_2_113, // sfix19_En18 
    input [18:0] Wgt_2_114, // sfix19_En18 
    input [18:0] Wgt_2_115, // sfix19_En18 
    input [18:0] Wgt_2_116, // sfix19_En18 
    input [18:0] Wgt_2_117, // sfix19_En18 
    input [18:0] Wgt_2_118, // sfix19_En18 
    input [18:0] Wgt_2_119, // sfix19_En18 
    input [18:0] Wgt_2_120, // sfix19_En18 
    input [18:0] Wgt_2_121, // sfix19_En18 
    input [18:0] Wgt_2_122, // sfix19_En18 
    input [18:0] Wgt_2_123, // sfix19_En18 
    input [18:0] Wgt_2_124, // sfix19_En18 
    input [18:0] Wgt_2_125, // sfix19_En18 
    input [18:0] Wgt_2_126, // sfix19_En18 
    input [18:0] Wgt_2_127, // sfix19_En18 
    input [18:0] Wgt_2_128, // sfix19_En18 
    input [18:0] Wgt_2_129, // sfix19_En18 
    input [18:0] Wgt_2_130, // sfix19_En18 
    input [18:0] Wgt_2_131, // sfix19_En18 
    input [18:0] Wgt_2_132, // sfix19_En18 
    input [18:0] Wgt_2_133, // sfix19_En18 
    input [18:0] Wgt_2_134, // sfix19_En18 
    input [18:0] Wgt_2_135, // sfix19_En18 
    input [18:0] Wgt_2_136, // sfix19_En18 
    input [18:0] Wgt_2_137, // sfix19_En18 
    input [18:0] Wgt_2_138, // sfix19_En18 
    input [18:0] Wgt_2_139, // sfix19_En18 
    input [18:0] Wgt_2_140, // sfix19_En18 
    input [18:0] Wgt_2_141, // sfix19_En18 
    input [18:0] Wgt_2_142, // sfix19_En18 
    input [18:0] Wgt_2_143, // sfix19_En18 
    input [18:0] Wgt_2_144, // sfix19_En18 
    input [18:0] Wgt_2_145, // sfix19_En18 
    input [18:0] Wgt_2_146, // sfix19_En18 
    input [18:0] Wgt_2_147, // sfix19_En18 
    input [18:0] Wgt_2_148, // sfix19_En18 
    input [18:0] Wgt_2_149, // sfix19_En18 
    input [18:0] Wgt_2_150, // sfix19_En18 
    input [18:0] Wgt_2_151, // sfix19_En18 
    input [18:0] Wgt_2_152, // sfix19_En18 
    input [18:0] Wgt_2_153, // sfix19_En18 
    input [18:0] Wgt_2_154, // sfix19_En18 
    input [18:0] Wgt_2_155, // sfix19_En18 
    input [18:0] Wgt_2_156, // sfix19_En18 
    input [18:0] Wgt_2_157, // sfix19_En18 
    input [18:0] Wgt_2_158, // sfix19_En18 
    input [18:0] Wgt_2_159, // sfix19_En18 
    input [18:0] Wgt_2_160, // sfix19_En18 
    input [18:0] Wgt_2_161, // sfix19_En18 
    input [18:0] Wgt_2_162, // sfix19_En18 
    input [18:0] Wgt_2_163, // sfix19_En18 
    input [18:0] Wgt_2_164, // sfix19_En18 
    input [18:0] Wgt_2_165, // sfix19_En18 
    input [18:0] Wgt_2_166, // sfix19_En18 
    input [18:0] Wgt_2_167, // sfix19_En18 
    input [18:0] Wgt_2_168, // sfix19_En18 
    input [18:0] Wgt_2_169, // sfix19_En18 
    input [18:0] Wgt_2_170, // sfix19_En18 
    input [18:0] Wgt_2_171, // sfix19_En18 
    input [18:0] Wgt_2_172, // sfix19_En18 
    input [18:0] Wgt_2_173, // sfix19_En18 
    input [18:0] Wgt_2_174, // sfix19_En18 
    input [18:0] Wgt_2_175, // sfix19_En18 
    input [18:0] Wgt_2_176, // sfix19_En18 
    input [18:0] Wgt_2_177, // sfix19_En18 
    input [18:0] Wgt_2_178, // sfix19_En18 
    input [18:0] Wgt_2_179, // sfix19_En18 
    input [18:0] Wgt_2_180, // sfix19_En18 
    input [18:0] Wgt_2_181, // sfix19_En18 
    input [18:0] Wgt_2_182, // sfix19_En18 
    input [18:0] Wgt_2_183, // sfix19_En18 
    input [18:0] Wgt_2_184, // sfix19_En18 
    input [18:0] Wgt_2_185, // sfix19_En18 
    input [18:0] Wgt_2_186, // sfix19_En18 
    input [18:0] Wgt_2_187, // sfix19_En18 
    input [18:0] Wgt_2_188, // sfix19_En18 
    input [18:0] Wgt_2_189, // sfix19_En18 
    input [18:0] Wgt_2_190, // sfix19_En18 
    input [18:0] Wgt_2_191, // sfix19_En18 
    input [18:0] Wgt_2_192, // sfix19_En18 
    input [18:0] Wgt_2_193, // sfix19_En18 
    input [18:0] Wgt_2_194, // sfix19_En18 
    input [18:0] Wgt_2_195, // sfix19_En18 
    input [18:0] Wgt_2_196, // sfix19_En18 
    input [18:0] Wgt_2_197, // sfix19_En18 
    input [18:0] Wgt_2_198, // sfix19_En18 
    input [18:0] Wgt_2_199, // sfix19_En18 
    input [18:0] Wgt_2_200, // sfix19_En18 
    input [18:0] Wgt_2_201, // sfix19_En18 
    input [18:0] Wgt_2_202, // sfix19_En18 
    input [18:0] Wgt_2_203, // sfix19_En18 
    input [18:0] Wgt_2_204, // sfix19_En18 
    input [18:0] Wgt_2_205, // sfix19_En18 
    input [18:0] Wgt_2_206, // sfix19_En18 
    input [18:0] Wgt_2_207, // sfix19_En18 
    input [18:0] Wgt_2_208, // sfix19_En18 
    input [18:0] Wgt_2_209, // sfix19_En18 
    input [18:0] Wgt_2_210, // sfix19_En18 
    input [18:0] Wgt_2_211, // sfix19_En18 
    input [18:0] Wgt_2_212, // sfix19_En18 
    input [18:0] Wgt_2_213, // sfix19_En18 
    input [18:0] Wgt_2_214, // sfix19_En18 
    input [18:0] Wgt_2_215, // sfix19_En18 
    input [18:0] Wgt_2_216, // sfix19_En18 
    input [18:0] Wgt_2_217, // sfix19_En18 
    input [18:0] Wgt_2_218, // sfix19_En18 
    input [18:0] Wgt_2_219, // sfix19_En18 
    input [18:0] Wgt_2_220, // sfix19_En18 
    input [18:0] Wgt_2_221, // sfix19_En18 
    input [18:0] Wgt_2_222, // sfix19_En18 
    input [18:0] Wgt_2_223, // sfix19_En18 
    input [18:0] Wgt_2_224, // sfix19_En18 
    input [18:0] Wgt_2_225, // sfix19_En18 
    input [18:0] Wgt_2_226, // sfix19_En18 
    input [18:0] Wgt_2_227, // sfix19_En18 
    input [18:0] Wgt_2_228, // sfix19_En18 
    input [18:0] Wgt_2_229, // sfix19_En18 
    input [18:0] Wgt_2_230, // sfix19_En18 
    input [18:0] Wgt_2_231, // sfix19_En18 
    input [18:0] Wgt_2_232, // sfix19_En18 
    input [18:0] Wgt_2_233, // sfix19_En18 
    input [18:0] Wgt_2_234, // sfix19_En18 
    input [18:0] Wgt_2_235, // sfix19_En18 
    input [18:0] Wgt_2_236, // sfix19_En18 
    input [18:0] Wgt_2_237, // sfix19_En18 
    input [18:0] Wgt_2_238, // sfix19_En18 
    input [18:0] Wgt_2_239, // sfix19_En18 
    input [18:0] Wgt_2_240, // sfix19_En18 
    input [18:0] Wgt_2_241, // sfix19_En18 
    input [18:0] Wgt_2_242, // sfix19_En18 
    input [18:0] Wgt_2_243, // sfix19_En18 
    input [18:0] Wgt_2_244, // sfix19_En18 
    input [18:0] Wgt_2_245, // sfix19_En18 
    input [18:0] Wgt_2_246, // sfix19_En18 
    input [18:0] Wgt_2_247, // sfix19_En18 
    input [18:0] Wgt_2_248, // sfix19_En18 
    input [18:0] Wgt_2_249, // sfix19_En18 
    input [18:0] Wgt_2_250, // sfix19_En18 
    input [18:0] Wgt_2_251, // sfix19_En18 
    input [18:0] Wgt_2_252, // sfix19_En18 
    input [18:0] Wgt_2_253, // sfix19_En18 
    input [18:0] Wgt_2_254, // sfix19_En18 
    input [18:0] Wgt_2_255, // sfix19_En18 
    input [18:0] Wgt_2_256, // sfix19_En18 
    input [18:0] Wgt_2_257, // sfix19_En18 
    input [18:0] Wgt_2_258, // sfix19_En18 
    input [18:0] Wgt_2_259, // sfix19_En18 
    input [18:0] Wgt_2_260, // sfix19_En18 
    input [18:0] Wgt_2_261, // sfix19_En18 
    input [18:0] Wgt_2_262, // sfix19_En18 
    input [18:0] Wgt_2_263, // sfix19_En18 
    input [18:0] Wgt_2_264, // sfix19_En18 
    input [18:0] Wgt_2_265, // sfix19_En18 
    input [18:0] Wgt_2_266, // sfix19_En18 
    input [18:0] Wgt_2_267, // sfix19_En18 
    input [18:0] Wgt_2_268, // sfix19_En18 
    input [18:0] Wgt_2_269, // sfix19_En18 
    input [18:0] Wgt_2_270, // sfix19_En18 
    input [18:0] Wgt_2_271, // sfix19_En18 
    input [18:0] Wgt_2_272, // sfix19_En18 
    input [18:0] Wgt_2_273, // sfix19_En18 
    input [18:0] Wgt_2_274, // sfix19_En18 
    input [18:0] Wgt_2_275, // sfix19_En18 
    input [18:0] Wgt_2_276, // sfix19_En18 
    input [18:0] Wgt_2_277, // sfix19_En18 
    input [18:0] Wgt_2_278, // sfix19_En18 
    input [18:0] Wgt_2_279, // sfix19_En18 
    input [18:0] Wgt_2_280, // sfix19_En18 
    input [18:0] Wgt_2_281, // sfix19_En18 
    input [18:0] Wgt_2_282, // sfix19_En18 
    input [18:0] Wgt_2_283, // sfix19_En18 
    input [18:0] Wgt_2_284, // sfix19_En18 
    input [18:0] Wgt_2_285, // sfix19_En18 
    input [18:0] Wgt_2_286, // sfix19_En18 
    input [18:0] Wgt_2_287, // sfix19_En18 
    input [18:0] Wgt_2_288, // sfix19_En18 
    input [18:0] Wgt_2_289, // sfix19_En18 
    input [18:0] Wgt_2_290, // sfix19_En18 
    input [18:0] Wgt_2_291, // sfix19_En18 
    input [18:0] Wgt_2_292, // sfix19_En18 
    input [18:0] Wgt_2_293, // sfix19_En18 
    input [18:0] Wgt_2_294, // sfix19_En18 
    input [18:0] Wgt_2_295, // sfix19_En18 
    input [18:0] Wgt_2_296, // sfix19_En18 
    input [18:0] Wgt_2_297, // sfix19_En18 
    input [18:0] Wgt_2_298, // sfix19_En18 
    input [18:0] Wgt_2_299, // sfix19_En18 
    input [18:0] Wgt_2_300, // sfix19_En18 
    input [18:0] Wgt_2_301, // sfix19_En18 
    input [18:0] Wgt_2_302, // sfix19_En18 
    input [18:0] Wgt_2_303, // sfix19_En18 
    input [18:0] Wgt_2_304, // sfix19_En18 
    input [18:0] Wgt_2_305, // sfix19_En18 
    input [18:0] Wgt_2_306, // sfix19_En18 
    input [18:0] Wgt_2_307, // sfix19_En18 
    input [18:0] Wgt_2_308, // sfix19_En18 
    input [18:0] Wgt_2_309, // sfix19_En18 
    input [18:0] Wgt_2_310, // sfix19_En18 
    input [18:0] Wgt_2_311, // sfix19_En18 
    input [18:0] Wgt_2_312, // sfix19_En18 
    input [18:0] Wgt_2_313, // sfix19_En18 
    input [18:0] Wgt_2_314, // sfix19_En18 
    input [18:0] Wgt_2_315, // sfix19_En18 
    input [18:0] Wgt_2_316, // sfix19_En18 
    input [18:0] Wgt_2_317, // sfix19_En18 
    input [18:0] Wgt_2_318, // sfix19_En18 
    input [18:0] Wgt_2_319, // sfix19_En18 
    input [18:0] Wgt_2_320, // sfix19_En18 
    input [18:0] Wgt_2_321, // sfix19_En18 
    input [18:0] Wgt_2_322, // sfix19_En18 
    input [18:0] Wgt_2_323, // sfix19_En18 
    input [18:0] Wgt_2_324, // sfix19_En18 
    input [18:0] Wgt_2_325, // sfix19_En18 
    input [18:0] Wgt_2_326, // sfix19_En18 
    input [18:0] Wgt_2_327, // sfix19_En18 
    input [18:0] Wgt_2_328, // sfix19_En18 
    input [18:0] Wgt_2_329, // sfix19_En18 
    input [18:0] Wgt_2_330, // sfix19_En18 
    input [18:0] Wgt_2_331, // sfix19_En18 
    input [18:0] Wgt_2_332, // sfix19_En18 
    input [18:0] Wgt_2_333, // sfix19_En18 
    input [18:0] Wgt_2_334, // sfix19_En18 
    input [18:0] Wgt_2_335, // sfix19_En18 
    input [18:0] Wgt_2_336, // sfix19_En18 
    input [18:0] Wgt_2_337, // sfix19_En18 
    input [18:0] Wgt_2_338, // sfix19_En18 
    input [18:0] Wgt_2_339, // sfix19_En18 
    input [18:0] Wgt_2_340, // sfix19_En18 
    input [18:0] Wgt_2_341, // sfix19_En18 
    input [18:0] Wgt_2_342, // sfix19_En18 
    input [18:0] Wgt_2_343, // sfix19_En18 
    input [18:0] Wgt_2_344, // sfix19_En18 
    input [18:0] Wgt_2_345, // sfix19_En18 
    input [18:0] Wgt_2_346, // sfix19_En18 
    input [18:0] Wgt_2_347, // sfix19_En18 
    input [18:0] Wgt_2_348, // sfix19_En18 
    input [18:0] Wgt_2_349, // sfix19_En18 
    input [18:0] Wgt_2_350, // sfix19_En18 
    input [18:0] Wgt_2_351, // sfix19_En18 
    input [18:0] Wgt_2_352, // sfix19_En18 
    input [18:0] Wgt_2_353, // sfix19_En18 
    input [18:0] Wgt_2_354, // sfix19_En18 
    input [18:0] Wgt_2_355, // sfix19_En18 
    input [18:0] Wgt_2_356, // sfix19_En18 
    input [18:0] Wgt_2_357, // sfix19_En18 
    input [18:0] Wgt_2_358, // sfix19_En18 
    input [18:0] Wgt_2_359, // sfix19_En18 
    input [18:0] Wgt_2_360, // sfix19_En18 
    input [18:0] Wgt_2_361, // sfix19_En18 
    input [18:0] Wgt_2_362, // sfix19_En18 
    input [18:0] Wgt_2_363, // sfix19_En18 
    input [18:0] Wgt_2_364, // sfix19_En18 
    input [18:0] Wgt_2_365, // sfix19_En18 
    input [18:0] Wgt_2_366, // sfix19_En18 
    input [18:0] Wgt_2_367, // sfix19_En18 
    input [18:0] Wgt_2_368, // sfix19_En18 
    input [18:0] Wgt_2_369, // sfix19_En18 
    input [18:0] Wgt_2_370, // sfix19_En18 
    input [18:0] Wgt_2_371, // sfix19_En18 
    input [18:0] Wgt_2_372, // sfix19_En18 
    input [18:0] Wgt_2_373, // sfix19_En18 
    input [18:0] Wgt_2_374, // sfix19_En18 
    input [18:0] Wgt_2_375, // sfix19_En18 
    input [18:0] Wgt_2_376, // sfix19_En18 
    input [18:0] Wgt_2_377, // sfix19_En18 
    input [18:0] Wgt_2_378, // sfix19_En18 
    input [18:0] Wgt_2_379, // sfix19_En18 
    input [18:0] Wgt_2_380, // sfix19_En18 
    input [18:0] Wgt_2_381, // sfix19_En18 
    input [18:0] Wgt_2_382, // sfix19_En18 
    input [18:0] Wgt_2_383, // sfix19_En18 
    input [18:0] Wgt_2_384, // sfix19_En18 
    input [18:0] Wgt_2_385, // sfix19_En18 
    input [18:0] Wgt_2_386, // sfix19_En18 
    input [18:0] Wgt_2_387, // sfix19_En18 
    input [18:0] Wgt_2_388, // sfix19_En18 
    input [18:0] Wgt_2_389, // sfix19_En18 
    input [18:0] Wgt_2_390, // sfix19_En18 
    input [18:0] Wgt_2_391, // sfix19_En18 
    input [18:0] Wgt_2_392, // sfix19_En18 
    input [18:0] Wgt_2_393, // sfix19_En18 
    input [18:0] Wgt_2_394, // sfix19_En18 
    input [18:0] Wgt_2_395, // sfix19_En18 
    input [18:0] Wgt_2_396, // sfix19_En18 
    input [18:0] Wgt_2_397, // sfix19_En18 
    input [18:0] Wgt_2_398, // sfix19_En18 
    input [18:0] Wgt_2_399, // sfix19_En18 
    input [18:0] Wgt_2_400, // sfix19_En18 
    input [18:0] Wgt_2_401, // sfix19_En18 
    input [18:0] Wgt_2_402, // sfix19_En18 
    input [18:0] Wgt_2_403, // sfix19_En18 
    input [18:0] Wgt_2_404, // sfix19_En18 
    input [18:0] Wgt_2_405, // sfix19_En18 
    input [18:0] Wgt_2_406, // sfix19_En18 
    input [18:0] Wgt_2_407, // sfix19_En18 
    input [18:0] Wgt_2_408, // sfix19_En18 
    input [18:0] Wgt_2_409, // sfix19_En18 
    input [18:0] Wgt_2_410, // sfix19_En18 
    input [18:0] Wgt_2_411, // sfix19_En18 
    input [18:0] Wgt_2_412, // sfix19_En18 
    input [18:0] Wgt_2_413, // sfix19_En18 
    input [18:0] Wgt_2_414, // sfix19_En18 
    input [18:0] Wgt_2_415, // sfix19_En18 
    input [18:0] Wgt_2_416, // sfix19_En18 
    input [18:0] Wgt_2_417, // sfix19_En18 
    input [18:0] Wgt_2_418, // sfix19_En18 
    input [18:0] Wgt_2_419, // sfix19_En18 
    input [18:0] Wgt_2_420, // sfix19_En18 
    input [18:0] Wgt_2_421, // sfix19_En18 
    input [18:0] Wgt_2_422, // sfix19_En18 
    input [18:0] Wgt_2_423, // sfix19_En18 
    input [18:0] Wgt_2_424, // sfix19_En18 
    input [18:0] Wgt_2_425, // sfix19_En18 
    input [18:0] Wgt_2_426, // sfix19_En18 
    input [18:0] Wgt_2_427, // sfix19_En18 
    input [18:0] Wgt_2_428, // sfix19_En18 
    input [18:0] Wgt_2_429, // sfix19_En18 
    input [18:0] Wgt_2_430, // sfix19_En18 
    input [18:0] Wgt_2_431, // sfix19_En18 
    input [18:0] Wgt_2_432, // sfix19_En18 
    input [18:0] Wgt_2_433, // sfix19_En18 
    input [18:0] Wgt_2_434, // sfix19_En18 
    input [18:0] Wgt_2_435, // sfix19_En18 
    input [18:0] Wgt_2_436, // sfix19_En18 
    input [18:0] Wgt_2_437, // sfix19_En18 
    input [18:0] Wgt_2_438, // sfix19_En18 
    input [18:0] Wgt_2_439, // sfix19_En18 
    input [18:0] Wgt_2_440, // sfix19_En18 
    input [18:0] Wgt_2_441, // sfix19_En18 
    input [18:0] Wgt_2_442, // sfix19_En18 
    input [18:0] Wgt_2_443, // sfix19_En18 
    input [18:0] Wgt_2_444, // sfix19_En18 
    input [18:0] Wgt_2_445, // sfix19_En18 
    input [18:0] Wgt_2_446, // sfix19_En18 
    input [18:0] Wgt_2_447, // sfix19_En18 
    input [18:0] Wgt_2_448, // sfix19_En18 
    input [18:0] Wgt_2_449, // sfix19_En18 
    input [18:0] Wgt_2_450, // sfix19_En18 
    input [18:0] Wgt_2_451, // sfix19_En18 
    input [18:0] Wgt_2_452, // sfix19_En18 
    input [18:0] Wgt_2_453, // sfix19_En18 
    input [18:0] Wgt_2_454, // sfix19_En18 
    input [18:0] Wgt_2_455, // sfix19_En18 
    input [18:0] Wgt_2_456, // sfix19_En18 
    input [18:0] Wgt_2_457, // sfix19_En18 
    input [18:0] Wgt_2_458, // sfix19_En18 
    input [18:0] Wgt_2_459, // sfix19_En18 
    input [18:0] Wgt_2_460, // sfix19_En18 
    input [18:0] Wgt_2_461, // sfix19_En18 
    input [18:0] Wgt_2_462, // sfix19_En18 
    input [18:0] Wgt_2_463, // sfix19_En18 
    input [18:0] Wgt_2_464, // sfix19_En18 
    input [18:0] Wgt_2_465, // sfix19_En18 
    input [18:0] Wgt_2_466, // sfix19_En18 
    input [18:0] Wgt_2_467, // sfix19_En18 
    input [18:0] Wgt_2_468, // sfix19_En18 
    input [18:0] Wgt_2_469, // sfix19_En18 
    input [18:0] Wgt_2_470, // sfix19_En18 
    input [18:0] Wgt_2_471, // sfix19_En18 
    input [18:0] Wgt_2_472, // sfix19_En18 
    input [18:0] Wgt_2_473, // sfix19_En18 
    input [18:0] Wgt_2_474, // sfix19_En18 
    input [18:0] Wgt_2_475, // sfix19_En18 
    input [18:0] Wgt_2_476, // sfix19_En18 
    input [18:0] Wgt_2_477, // sfix19_En18 
    input [18:0] Wgt_2_478, // sfix19_En18 
    input [18:0] Wgt_2_479, // sfix19_En18 
    input [18:0] Wgt_2_480, // sfix19_En18 
    input [18:0] Wgt_2_481, // sfix19_En18 
    input [18:0] Wgt_2_482, // sfix19_En18 
    input [18:0] Wgt_2_483, // sfix19_En18 
    input [18:0] Wgt_2_484, // sfix19_En18 
    input [18:0] Wgt_2_485, // sfix19_En18 
    input [18:0] Wgt_2_486, // sfix19_En18 
    input [18:0] Wgt_2_487, // sfix19_En18 
    input [18:0] Wgt_2_488, // sfix19_En18 
    input [18:0] Wgt_2_489, // sfix19_En18 
    input [18:0] Wgt_2_490, // sfix19_En18 
    input [18:0] Wgt_2_491, // sfix19_En18 
    input [18:0] Wgt_2_492, // sfix19_En18 
    input [18:0] Wgt_2_493, // sfix19_En18 
    input [18:0] Wgt_2_494, // sfix19_En18 
    input [18:0] Wgt_2_495, // sfix19_En18 
    input [18:0] Wgt_2_496, // sfix19_En18 
    input [18:0] Wgt_2_497, // sfix19_En18 
    input [18:0] Wgt_2_498, // sfix19_En18 
    input [18:0] Wgt_2_499, // sfix19_En18 
    input [18:0] Wgt_2_500, // sfix19_En18 
    input [18:0] Wgt_2_501, // sfix19_En18 
    input [18:0] Wgt_2_502, // sfix19_En18 
    input [18:0] Wgt_2_503, // sfix19_En18 
    input [18:0] Wgt_2_504, // sfix19_En18 
    input [18:0] Wgt_2_505, // sfix19_En18 
    input [18:0] Wgt_2_506, // sfix19_En18 
    input [18:0] Wgt_2_507, // sfix19_En18 
    input [18:0] Wgt_2_508, // sfix19_En18 
    input [18:0] Wgt_2_509, // sfix19_En18 
    input [18:0] Wgt_2_510, // sfix19_En18 
    input [18:0] Wgt_2_511, // sfix19_En18 
    input [18:0] Wgt_2_512, // sfix19_En18 
    input [18:0] Wgt_2_513, // sfix19_En18 
    input [18:0] Wgt_2_514, // sfix19_En18 
    input [18:0] Wgt_2_515, // sfix19_En18 
    input [18:0] Wgt_2_516, // sfix19_En18 
    input [18:0] Wgt_2_517, // sfix19_En18 
    input [18:0] Wgt_2_518, // sfix19_En18 
    input [18:0] Wgt_2_519, // sfix19_En18 
    input [18:0] Wgt_2_520, // sfix19_En18 
    input [18:0] Wgt_2_521, // sfix19_En18 
    input [18:0] Wgt_2_522, // sfix19_En18 
    input [18:0] Wgt_2_523, // sfix19_En18 
    input [18:0] Wgt_2_524, // sfix19_En18 
    input [18:0] Wgt_2_525, // sfix19_En18 
    input [18:0] Wgt_2_526, // sfix19_En18 
    input [18:0] Wgt_2_527, // sfix19_En18 
    input [18:0] Wgt_2_528, // sfix19_En18 
    input [18:0] Wgt_2_529, // sfix19_En18 
    input [18:0] Wgt_2_530, // sfix19_En18 
    input [18:0] Wgt_2_531, // sfix19_En18 
    input [18:0] Wgt_2_532, // sfix19_En18 
    input [18:0] Wgt_2_533, // sfix19_En18 
    input [18:0] Wgt_2_534, // sfix19_En18 
    input [18:0] Wgt_2_535, // sfix19_En18 
    input [18:0] Wgt_2_536, // sfix19_En18 
    input [18:0] Wgt_2_537, // sfix19_En18 
    input [18:0] Wgt_2_538, // sfix19_En18 
    input [18:0] Wgt_2_539, // sfix19_En18 
    input [18:0] Wgt_2_540, // sfix19_En18 
    input [18:0] Wgt_2_541, // sfix19_En18 
    input [18:0] Wgt_2_542, // sfix19_En18 
    input [18:0] Wgt_2_543, // sfix19_En18 
    input [18:0] Wgt_2_544, // sfix19_En18 
    input [18:0] Wgt_2_545, // sfix19_En18 
    input [18:0] Wgt_2_546, // sfix19_En18 
    input [18:0] Wgt_2_547, // sfix19_En18 
    input [18:0] Wgt_2_548, // sfix19_En18 
    input [18:0] Wgt_2_549, // sfix19_En18 
    input [18:0] Wgt_2_550, // sfix19_En18 
    input [18:0] Wgt_2_551, // sfix19_En18 
    input [18:0] Wgt_2_552, // sfix19_En18 
    input [18:0] Wgt_2_553, // sfix19_En18 
    input [18:0] Wgt_2_554, // sfix19_En18 
    input [18:0] Wgt_2_555, // sfix19_En18 
    input [18:0] Wgt_2_556, // sfix19_En18 
    input [18:0] Wgt_2_557, // sfix19_En18 
    input [18:0] Wgt_2_558, // sfix19_En18 
    input [18:0] Wgt_2_559, // sfix19_En18 
    input [18:0] Wgt_2_560, // sfix19_En18 
    input [18:0] Wgt_2_561, // sfix19_En18 
    input [18:0] Wgt_2_562, // sfix19_En18 
    input [18:0] Wgt_2_563, // sfix19_En18 
    input [18:0] Wgt_2_564, // sfix19_En18 
    input [18:0] Wgt_2_565, // sfix19_En18 
    input [18:0] Wgt_2_566, // sfix19_En18 
    input [18:0] Wgt_2_567, // sfix19_En18 
    input [18:0] Wgt_2_568, // sfix19_En18 
    input [18:0] Wgt_2_569, // sfix19_En18 
    input [18:0] Wgt_2_570, // sfix19_En18 
    input [18:0] Wgt_2_571, // sfix19_En18 
    input [18:0] Wgt_2_572, // sfix19_En18 
    input [18:0] Wgt_2_573, // sfix19_En18 
    input [18:0] Wgt_2_574, // sfix19_En18 
    input [18:0] Wgt_2_575, // sfix19_En18 
    input [18:0] Wgt_2_576, // sfix19_En18 
    input [18:0] Wgt_2_577, // sfix19_En18 
    input [18:0] Wgt_2_578, // sfix19_En18 
    input [18:0] Wgt_2_579, // sfix19_En18 
    input [18:0] Wgt_2_580, // sfix19_En18 
    input [18:0] Wgt_2_581, // sfix19_En18 
    input [18:0] Wgt_2_582, // sfix19_En18 
    input [18:0] Wgt_2_583, // sfix19_En18 
    input [18:0] Wgt_2_584, // sfix19_En18 
    input [18:0] Wgt_2_585, // sfix19_En18 
    input [18:0] Wgt_2_586, // sfix19_En18 
    input [18:0] Wgt_2_587, // sfix19_En18 
    input [18:0] Wgt_2_588, // sfix19_En18 
    input [18:0] Wgt_2_589, // sfix19_En18 
    input [18:0] Wgt_2_590, // sfix19_En18 
    input [18:0] Wgt_2_591, // sfix19_En18 
    input [18:0] Wgt_2_592, // sfix19_En18 
    input [18:0] Wgt_2_593, // sfix19_En18 
    input [18:0] Wgt_2_594, // sfix19_En18 
    input [18:0] Wgt_2_595, // sfix19_En18 
    input [18:0] Wgt_2_596, // sfix19_En18 
    input [18:0] Wgt_2_597, // sfix19_En18 
    input [18:0] Wgt_2_598, // sfix19_En18 
    input [18:0] Wgt_2_599, // sfix19_En18 
    input [18:0] Wgt_2_600, // sfix19_En18 
    input [18:0] Wgt_2_601, // sfix19_En18 
    input [18:0] Wgt_2_602, // sfix19_En18 
    input [18:0] Wgt_2_603, // sfix19_En18 
    input [18:0] Wgt_2_604, // sfix19_En18 
    input [18:0] Wgt_2_605, // sfix19_En18 
    input [18:0] Wgt_2_606, // sfix19_En18 
    input [18:0] Wgt_2_607, // sfix19_En18 
    input [18:0] Wgt_2_608, // sfix19_En18 
    input [18:0] Wgt_2_609, // sfix19_En18 
    input [18:0] Wgt_2_610, // sfix19_En18 
    input [18:0] Wgt_2_611, // sfix19_En18 
    input [18:0] Wgt_2_612, // sfix19_En18 
    input [18:0] Wgt_2_613, // sfix19_En18 
    input [18:0] Wgt_2_614, // sfix19_En18 
    input [18:0] Wgt_2_615, // sfix19_En18 
    input [18:0] Wgt_2_616, // sfix19_En18 
    input [18:0] Wgt_2_617, // sfix19_En18 
    input [18:0] Wgt_2_618, // sfix19_En18 
    input [18:0] Wgt_2_619, // sfix19_En18 
    input [18:0] Wgt_2_620, // sfix19_En18 
    input [18:0] Wgt_2_621, // sfix19_En18 
    input [18:0] Wgt_2_622, // sfix19_En18 
    input [18:0] Wgt_2_623, // sfix19_En18 
    input [18:0] Wgt_2_624, // sfix19_En18 
    input [18:0] Wgt_2_625, // sfix19_En18 
    input [18:0] Wgt_2_626, // sfix19_En18 
    input [18:0] Wgt_2_627, // sfix19_En18 
    input [18:0] Wgt_2_628, // sfix19_En18 
    input [18:0] Wgt_2_629, // sfix19_En18 
    input [18:0] Wgt_2_630, // sfix19_En18 
    input [18:0] Wgt_2_631, // sfix19_En18 
    input [18:0] Wgt_2_632, // sfix19_En18 
    input [18:0] Wgt_2_633, // sfix19_En18 
    input [18:0] Wgt_2_634, // sfix19_En18 
    input [18:0] Wgt_2_635, // sfix19_En18 
    input [18:0] Wgt_2_636, // sfix19_En18 
    input [18:0] Wgt_2_637, // sfix19_En18 
    input [18:0] Wgt_2_638, // sfix19_En18 
    input [18:0] Wgt_2_639, // sfix19_En18 
    input [18:0] Wgt_2_640, // sfix19_En18 
    input [18:0] Wgt_2_641, // sfix19_En18 
    input [18:0] Wgt_2_642, // sfix19_En18 
    input [18:0] Wgt_2_643, // sfix19_En18 
    input [18:0] Wgt_2_644, // sfix19_En18 
    input [18:0] Wgt_2_645, // sfix19_En18 
    input [18:0] Wgt_2_646, // sfix19_En18 
    input [18:0] Wgt_2_647, // sfix19_En18 
    input [18:0] Wgt_2_648, // sfix19_En18 
    input [18:0] Wgt_2_649, // sfix19_En18 
    input [18:0] Wgt_2_650, // sfix19_En18 
    input [18:0] Wgt_2_651, // sfix19_En18 
    input [18:0] Wgt_2_652, // sfix19_En18 
    input [18:0] Wgt_2_653, // sfix19_En18 
    input [18:0] Wgt_2_654, // sfix19_En18 
    input [18:0] Wgt_2_655, // sfix19_En18 
    input [18:0] Wgt_2_656, // sfix19_En18 
    input [18:0] Wgt_2_657, // sfix19_En18 
    input [18:0] Wgt_2_658, // sfix19_En18 
    input [18:0] Wgt_2_659, // sfix19_En18 
    input [18:0] Wgt_2_660, // sfix19_En18 
    input [18:0] Wgt_2_661, // sfix19_En18 
    input [18:0] Wgt_2_662, // sfix19_En18 
    input [18:0] Wgt_2_663, // sfix19_En18 
    input [18:0] Wgt_2_664, // sfix19_En18 
    input [18:0] Wgt_2_665, // sfix19_En18 
    input [18:0] Wgt_2_666, // sfix19_En18 
    input [18:0] Wgt_2_667, // sfix19_En18 
    input [18:0] Wgt_2_668, // sfix19_En18 
    input [18:0] Wgt_2_669, // sfix19_En18 
    input [18:0] Wgt_2_670, // sfix19_En18 
    input [18:0] Wgt_2_671, // sfix19_En18 
    input [18:0] Wgt_2_672, // sfix19_En18 
    input [18:0] Wgt_2_673, // sfix19_En18 
    input [18:0] Wgt_2_674, // sfix19_En18 
    input [18:0] Wgt_2_675, // sfix19_En18 
    input [18:0] Wgt_2_676, // sfix19_En18 
    input [18:0] Wgt_2_677, // sfix19_En18 
    input [18:0] Wgt_2_678, // sfix19_En18 
    input [18:0] Wgt_2_679, // sfix19_En18 
    input [18:0] Wgt_2_680, // sfix19_En18 
    input [18:0] Wgt_2_681, // sfix19_En18 
    input [18:0] Wgt_2_682, // sfix19_En18 
    input [18:0] Wgt_2_683, // sfix19_En18 
    input [18:0] Wgt_2_684, // sfix19_En18 
    input [18:0] Wgt_2_685, // sfix19_En18 
    input [18:0] Wgt_2_686, // sfix19_En18 
    input [18:0] Wgt_2_687, // sfix19_En18 
    input [18:0] Wgt_2_688, // sfix19_En18 
    input [18:0] Wgt_2_689, // sfix19_En18 
    input [18:0] Wgt_2_690, // sfix19_En18 
    input [18:0] Wgt_2_691, // sfix19_En18 
    input [18:0] Wgt_2_692, // sfix19_En18 
    input [18:0] Wgt_2_693, // sfix19_En18 
    input [18:0] Wgt_2_694, // sfix19_En18 
    input [18:0] Wgt_2_695, // sfix19_En18 
    input [18:0] Wgt_2_696, // sfix19_En18 
    input [18:0] Wgt_2_697, // sfix19_En18 
    input [18:0] Wgt_2_698, // sfix19_En18 
    input [18:0] Wgt_2_699, // sfix19_En18 
    input [18:0] Wgt_2_700, // sfix19_En18 
    input [18:0] Wgt_2_701, // sfix19_En18 
    input [18:0] Wgt_2_702, // sfix19_En18 
    input [18:0] Wgt_2_703, // sfix19_En18 
    input [18:0] Wgt_2_704, // sfix19_En18 
    input [18:0] Wgt_2_705, // sfix19_En18 
    input [18:0] Wgt_2_706, // sfix19_En18 
    input [18:0] Wgt_2_707, // sfix19_En18 
    input [18:0] Wgt_2_708, // sfix19_En18 
    input [18:0] Wgt_2_709, // sfix19_En18 
    input [18:0] Wgt_2_710, // sfix19_En18 
    input [18:0] Wgt_2_711, // sfix19_En18 
    input [18:0] Wgt_2_712, // sfix19_En18 
    input [18:0] Wgt_2_713, // sfix19_En18 
    input [18:0] Wgt_2_714, // sfix19_En18 
    input [18:0] Wgt_2_715, // sfix19_En18 
    input [18:0] Wgt_2_716, // sfix19_En18 
    input [18:0] Wgt_2_717, // sfix19_En18 
    input [18:0] Wgt_2_718, // sfix19_En18 
    input [18:0] Wgt_2_719, // sfix19_En18 
    input [18:0] Wgt_2_720, // sfix19_En18 
    input [18:0] Wgt_2_721, // sfix19_En18 
    input [18:0] Wgt_2_722, // sfix19_En18 
    input [18:0] Wgt_2_723, // sfix19_En18 
    input [18:0] Wgt_2_724, // sfix19_En18 
    input [18:0] Wgt_2_725, // sfix19_En18 
    input [18:0] Wgt_2_726, // sfix19_En18 
    input [18:0] Wgt_2_727, // sfix19_En18 
    input [18:0] Wgt_2_728, // sfix19_En18 
    input [18:0] Wgt_2_729, // sfix19_En18 
    input [18:0] Wgt_2_730, // sfix19_En18 
    input [18:0] Wgt_2_731, // sfix19_En18 
    input [18:0] Wgt_2_732, // sfix19_En18 
    input [18:0] Wgt_2_733, // sfix19_En18 
    input [18:0] Wgt_2_734, // sfix19_En18 
    input [18:0] Wgt_2_735, // sfix19_En18 
    input [18:0] Wgt_2_736, // sfix19_En18 
    input [18:0] Wgt_2_737, // sfix19_En18 
    input [18:0] Wgt_2_738, // sfix19_En18 
    input [18:0] Wgt_2_739, // sfix19_En18 
    input [18:0] Wgt_2_740, // sfix19_En18 
    input [18:0] Wgt_2_741, // sfix19_En18 
    input [18:0] Wgt_2_742, // sfix19_En18 
    input [18:0] Wgt_2_743, // sfix19_En18 
    input [18:0] Wgt_2_744, // sfix19_En18 
    input [18:0] Wgt_2_745, // sfix19_En18 
    input [18:0] Wgt_2_746, // sfix19_En18 
    input [18:0] Wgt_2_747, // sfix19_En18 
    input [18:0] Wgt_2_748, // sfix19_En18 
    input [18:0] Wgt_2_749, // sfix19_En18 
    input [18:0] Wgt_2_750, // sfix19_En18 
    input [18:0] Wgt_2_751, // sfix19_En18 
    input [18:0] Wgt_2_752, // sfix19_En18 
    input [18:0] Wgt_2_753, // sfix19_En18 
    input [18:0] Wgt_2_754, // sfix19_En18 
    input [18:0] Wgt_2_755, // sfix19_En18 
    input [18:0] Wgt_2_756, // sfix19_En18 
    input [18:0] Wgt_2_757, // sfix19_En18 
    input [18:0] Wgt_2_758, // sfix19_En18 
    input [18:0] Wgt_2_759, // sfix19_En18 
    input [18:0] Wgt_2_760, // sfix19_En18 
    input [18:0] Wgt_2_761, // sfix19_En18 
    input [18:0] Wgt_2_762, // sfix19_En18 
    input [18:0] Wgt_2_763, // sfix19_En18 
    input [18:0] Wgt_2_764, // sfix19_En18 
    input [18:0] Wgt_2_765, // sfix19_En18 
    input [18:0] Wgt_2_766, // sfix19_En18 
    input [18:0] Wgt_2_767, // sfix19_En18 
    input [18:0] Wgt_2_768, // sfix19_En18 
    input [18:0] Wgt_2_769, // sfix19_En18 
    input [18:0] Wgt_2_770, // sfix19_En18 
    input [18:0] Wgt_2_771, // sfix19_En18 
    input [18:0] Wgt_2_772, // sfix19_En18 
    input [18:0] Wgt_2_773, // sfix19_En18 
    input [18:0] Wgt_2_774, // sfix19_En18 
    input [18:0] Wgt_2_775, // sfix19_En18 
    input [18:0] Wgt_2_776, // sfix19_En18 
    input [18:0] Wgt_2_777, // sfix19_En18 
    input [18:0] Wgt_2_778, // sfix19_En18 
    input [18:0] Wgt_2_779, // sfix19_En18 
    input [18:0] Wgt_2_780, // sfix19_En18 
    input [18:0] Wgt_2_781, // sfix19_En18 
    input [18:0] Wgt_2_782, // sfix19_En18 
    input [18:0] Wgt_2_783, // sfix19_En18 
    input [18:0] Wgt_2_784, // sfix19_En18 
    input [18:0] Wgt_3_0, // sfix19_En18 
    input [18:0] Wgt_3_1, // sfix19_En18 
    input [18:0] Wgt_3_2, // sfix19_En18 
    input [18:0] Wgt_3_3, // sfix19_En18 
    input [18:0] Wgt_3_4, // sfix19_En18 
    input [18:0] Wgt_3_5, // sfix19_En18 
    input [18:0] Wgt_3_6, // sfix19_En18 
    input [18:0] Wgt_3_7, // sfix19_En18 
    input [18:0] Wgt_3_8, // sfix19_En18 
    input [18:0] Wgt_3_9, // sfix19_En18 
    input [18:0] Wgt_3_10, // sfix19_En18 
    input [18:0] Wgt_3_11, // sfix19_En18 
    input [18:0] Wgt_3_12, // sfix19_En18 
    input [18:0] Wgt_3_13, // sfix19_En18 
    input [18:0] Wgt_3_14, // sfix19_En18 
    input [18:0] Wgt_3_15, // sfix19_En18 
    input [18:0] Wgt_3_16, // sfix19_En18 
    input [18:0] Wgt_3_17, // sfix19_En18 
    input [18:0] Wgt_3_18, // sfix19_En18 
    input [18:0] Wgt_3_19, // sfix19_En18 
    input [18:0] Wgt_3_20, // sfix19_En18 
    input [18:0] Wgt_3_21, // sfix19_En18 
    input [18:0] Wgt_3_22, // sfix19_En18 
    input [18:0] Wgt_3_23, // sfix19_En18 
    input [18:0] Wgt_3_24, // sfix19_En18 
    input [18:0] Wgt_3_25, // sfix19_En18 
    input [18:0] Wgt_3_26, // sfix19_En18 
    input [18:0] Wgt_3_27, // sfix19_En18 
    input [18:0] Wgt_3_28, // sfix19_En18 
    input [18:0] Wgt_3_29, // sfix19_En18 
    input [18:0] Wgt_3_30, // sfix19_En18 
    input [18:0] Wgt_3_31, // sfix19_En18 
    input [18:0] Wgt_3_32, // sfix19_En18 
    input [18:0] Wgt_3_33, // sfix19_En18 
    input [18:0] Wgt_3_34, // sfix19_En18 
    input [18:0] Wgt_3_35, // sfix19_En18 
    input [18:0] Wgt_3_36, // sfix19_En18 
    input [18:0] Wgt_3_37, // sfix19_En18 
    input [18:0] Wgt_3_38, // sfix19_En18 
    input [18:0] Wgt_3_39, // sfix19_En18 
    input [18:0] Wgt_3_40, // sfix19_En18 
    input [18:0] Wgt_3_41, // sfix19_En18 
    input [18:0] Wgt_3_42, // sfix19_En18 
    input [18:0] Wgt_3_43, // sfix19_En18 
    input [18:0] Wgt_3_44, // sfix19_En18 
    input [18:0] Wgt_3_45, // sfix19_En18 
    input [18:0] Wgt_3_46, // sfix19_En18 
    input [18:0] Wgt_3_47, // sfix19_En18 
    input [18:0] Wgt_3_48, // sfix19_En18 
    input [18:0] Wgt_3_49, // sfix19_En18 
    input [18:0] Wgt_3_50, // sfix19_En18 
    input [18:0] Wgt_3_51, // sfix19_En18 
    input [18:0] Wgt_3_52, // sfix19_En18 
    input [18:0] Wgt_3_53, // sfix19_En18 
    input [18:0] Wgt_3_54, // sfix19_En18 
    input [18:0] Wgt_3_55, // sfix19_En18 
    input [18:0] Wgt_3_56, // sfix19_En18 
    input [18:0] Wgt_3_57, // sfix19_En18 
    input [18:0] Wgt_3_58, // sfix19_En18 
    input [18:0] Wgt_3_59, // sfix19_En18 
    input [18:0] Wgt_3_60, // sfix19_En18 
    input [18:0] Wgt_3_61, // sfix19_En18 
    input [18:0] Wgt_3_62, // sfix19_En18 
    input [18:0] Wgt_3_63, // sfix19_En18 
    input [18:0] Wgt_3_64, // sfix19_En18 
    input [18:0] Wgt_3_65, // sfix19_En18 
    input [18:0] Wgt_3_66, // sfix19_En18 
    input [18:0] Wgt_3_67, // sfix19_En18 
    input [18:0] Wgt_3_68, // sfix19_En18 
    input [18:0] Wgt_3_69, // sfix19_En18 
    input [18:0] Wgt_3_70, // sfix19_En18 
    input [18:0] Wgt_3_71, // sfix19_En18 
    input [18:0] Wgt_3_72, // sfix19_En18 
    input [18:0] Wgt_3_73, // sfix19_En18 
    input [18:0] Wgt_3_74, // sfix19_En18 
    input [18:0] Wgt_3_75, // sfix19_En18 
    input [18:0] Wgt_3_76, // sfix19_En18 
    input [18:0] Wgt_3_77, // sfix19_En18 
    input [18:0] Wgt_3_78, // sfix19_En18 
    input [18:0] Wgt_3_79, // sfix19_En18 
    input [18:0] Wgt_3_80, // sfix19_En18 
    input [18:0] Wgt_3_81, // sfix19_En18 
    input [18:0] Wgt_3_82, // sfix19_En18 
    input [18:0] Wgt_3_83, // sfix19_En18 
    input [18:0] Wgt_3_84, // sfix19_En18 
    input [18:0] Wgt_3_85, // sfix19_En18 
    input [18:0] Wgt_3_86, // sfix19_En18 
    input [18:0] Wgt_3_87, // sfix19_En18 
    input [18:0] Wgt_3_88, // sfix19_En18 
    input [18:0] Wgt_3_89, // sfix19_En18 
    input [18:0] Wgt_3_90, // sfix19_En18 
    input [18:0] Wgt_3_91, // sfix19_En18 
    input [18:0] Wgt_3_92, // sfix19_En18 
    input [18:0] Wgt_3_93, // sfix19_En18 
    input [18:0] Wgt_3_94, // sfix19_En18 
    input [18:0] Wgt_3_95, // sfix19_En18 
    input [18:0] Wgt_3_96, // sfix19_En18 
    input [18:0] Wgt_3_97, // sfix19_En18 
    input [18:0] Wgt_3_98, // sfix19_En18 
    input [18:0] Wgt_3_99, // sfix19_En18 
    input [18:0] Wgt_3_100, // sfix19_En18 
    input [18:0] Wgt_3_101, // sfix19_En18 
    input [18:0] Wgt_3_102, // sfix19_En18 
    input [18:0] Wgt_3_103, // sfix19_En18 
    input [18:0] Wgt_3_104, // sfix19_En18 
    input [18:0] Wgt_3_105, // sfix19_En18 
    input [18:0] Wgt_3_106, // sfix19_En18 
    input [18:0] Wgt_3_107, // sfix19_En18 
    input [18:0] Wgt_3_108, // sfix19_En18 
    input [18:0] Wgt_3_109, // sfix19_En18 
    input [18:0] Wgt_3_110, // sfix19_En18 
    input [18:0] Wgt_3_111, // sfix19_En18 
    input [18:0] Wgt_3_112, // sfix19_En18 
    input [18:0] Wgt_3_113, // sfix19_En18 
    input [18:0] Wgt_3_114, // sfix19_En18 
    input [18:0] Wgt_3_115, // sfix19_En18 
    input [18:0] Wgt_3_116, // sfix19_En18 
    input [18:0] Wgt_3_117, // sfix19_En18 
    input [18:0] Wgt_3_118, // sfix19_En18 
    input [18:0] Wgt_3_119, // sfix19_En18 
    input [18:0] Wgt_3_120, // sfix19_En18 
    input [18:0] Wgt_3_121, // sfix19_En18 
    input [18:0] Wgt_3_122, // sfix19_En18 
    input [18:0] Wgt_3_123, // sfix19_En18 
    input [18:0] Wgt_3_124, // sfix19_En18 
    input [18:0] Wgt_3_125, // sfix19_En18 
    input [18:0] Wgt_3_126, // sfix19_En18 
    input [18:0] Wgt_3_127, // sfix19_En18 
    input [18:0] Wgt_3_128, // sfix19_En18 
    input [18:0] Wgt_3_129, // sfix19_En18 
    input [18:0] Wgt_3_130, // sfix19_En18 
    input [18:0] Wgt_3_131, // sfix19_En18 
    input [18:0] Wgt_3_132, // sfix19_En18 
    input [18:0] Wgt_3_133, // sfix19_En18 
    input [18:0] Wgt_3_134, // sfix19_En18 
    input [18:0] Wgt_3_135, // sfix19_En18 
    input [18:0] Wgt_3_136, // sfix19_En18 
    input [18:0] Wgt_3_137, // sfix19_En18 
    input [18:0] Wgt_3_138, // sfix19_En18 
    input [18:0] Wgt_3_139, // sfix19_En18 
    input [18:0] Wgt_3_140, // sfix19_En18 
    input [18:0] Wgt_3_141, // sfix19_En18 
    input [18:0] Wgt_3_142, // sfix19_En18 
    input [18:0] Wgt_3_143, // sfix19_En18 
    input [18:0] Wgt_3_144, // sfix19_En18 
    input [18:0] Wgt_3_145, // sfix19_En18 
    input [18:0] Wgt_3_146, // sfix19_En18 
    input [18:0] Wgt_3_147, // sfix19_En18 
    input [18:0] Wgt_3_148, // sfix19_En18 
    input [18:0] Wgt_3_149, // sfix19_En18 
    input [18:0] Wgt_3_150, // sfix19_En18 
    input [18:0] Wgt_3_151, // sfix19_En18 
    input [18:0] Wgt_3_152, // sfix19_En18 
    input [18:0] Wgt_3_153, // sfix19_En18 
    input [18:0] Wgt_3_154, // sfix19_En18 
    input [18:0] Wgt_3_155, // sfix19_En18 
    input [18:0] Wgt_3_156, // sfix19_En18 
    input [18:0] Wgt_3_157, // sfix19_En18 
    input [18:0] Wgt_3_158, // sfix19_En18 
    input [18:0] Wgt_3_159, // sfix19_En18 
    input [18:0] Wgt_3_160, // sfix19_En18 
    input [18:0] Wgt_3_161, // sfix19_En18 
    input [18:0] Wgt_3_162, // sfix19_En18 
    input [18:0] Wgt_3_163, // sfix19_En18 
    input [18:0] Wgt_3_164, // sfix19_En18 
    input [18:0] Wgt_3_165, // sfix19_En18 
    input [18:0] Wgt_3_166, // sfix19_En18 
    input [18:0] Wgt_3_167, // sfix19_En18 
    input [18:0] Wgt_3_168, // sfix19_En18 
    input [18:0] Wgt_3_169, // sfix19_En18 
    input [18:0] Wgt_3_170, // sfix19_En18 
    input [18:0] Wgt_3_171, // sfix19_En18 
    input [18:0] Wgt_3_172, // sfix19_En18 
    input [18:0] Wgt_3_173, // sfix19_En18 
    input [18:0] Wgt_3_174, // sfix19_En18 
    input [18:0] Wgt_3_175, // sfix19_En18 
    input [18:0] Wgt_3_176, // sfix19_En18 
    input [18:0] Wgt_3_177, // sfix19_En18 
    input [18:0] Wgt_3_178, // sfix19_En18 
    input [18:0] Wgt_3_179, // sfix19_En18 
    input [18:0] Wgt_3_180, // sfix19_En18 
    input [18:0] Wgt_3_181, // sfix19_En18 
    input [18:0] Wgt_3_182, // sfix19_En18 
    input [18:0] Wgt_3_183, // sfix19_En18 
    input [18:0] Wgt_3_184, // sfix19_En18 
    input [18:0] Wgt_3_185, // sfix19_En18 
    input [18:0] Wgt_3_186, // sfix19_En18 
    input [18:0] Wgt_3_187, // sfix19_En18 
    input [18:0] Wgt_3_188, // sfix19_En18 
    input [18:0] Wgt_3_189, // sfix19_En18 
    input [18:0] Wgt_3_190, // sfix19_En18 
    input [18:0] Wgt_3_191, // sfix19_En18 
    input [18:0] Wgt_3_192, // sfix19_En18 
    input [18:0] Wgt_3_193, // sfix19_En18 
    input [18:0] Wgt_3_194, // sfix19_En18 
    input [18:0] Wgt_3_195, // sfix19_En18 
    input [18:0] Wgt_3_196, // sfix19_En18 
    input [18:0] Wgt_3_197, // sfix19_En18 
    input [18:0] Wgt_3_198, // sfix19_En18 
    input [18:0] Wgt_3_199, // sfix19_En18 
    input [18:0] Wgt_3_200, // sfix19_En18 
    input [18:0] Wgt_3_201, // sfix19_En18 
    input [18:0] Wgt_3_202, // sfix19_En18 
    input [18:0] Wgt_3_203, // sfix19_En18 
    input [18:0] Wgt_3_204, // sfix19_En18 
    input [18:0] Wgt_3_205, // sfix19_En18 
    input [18:0] Wgt_3_206, // sfix19_En18 
    input [18:0] Wgt_3_207, // sfix19_En18 
    input [18:0] Wgt_3_208, // sfix19_En18 
    input [18:0] Wgt_3_209, // sfix19_En18 
    input [18:0] Wgt_3_210, // sfix19_En18 
    input [18:0] Wgt_3_211, // sfix19_En18 
    input [18:0] Wgt_3_212, // sfix19_En18 
    input [18:0] Wgt_3_213, // sfix19_En18 
    input [18:0] Wgt_3_214, // sfix19_En18 
    input [18:0] Wgt_3_215, // sfix19_En18 
    input [18:0] Wgt_3_216, // sfix19_En18 
    input [18:0] Wgt_3_217, // sfix19_En18 
    input [18:0] Wgt_3_218, // sfix19_En18 
    input [18:0] Wgt_3_219, // sfix19_En18 
    input [18:0] Wgt_3_220, // sfix19_En18 
    input [18:0] Wgt_3_221, // sfix19_En18 
    input [18:0] Wgt_3_222, // sfix19_En18 
    input [18:0] Wgt_3_223, // sfix19_En18 
    input [18:0] Wgt_3_224, // sfix19_En18 
    input [18:0] Wgt_3_225, // sfix19_En18 
    input [18:0] Wgt_3_226, // sfix19_En18 
    input [18:0] Wgt_3_227, // sfix19_En18 
    input [18:0] Wgt_3_228, // sfix19_En18 
    input [18:0] Wgt_3_229, // sfix19_En18 
    input [18:0] Wgt_3_230, // sfix19_En18 
    input [18:0] Wgt_3_231, // sfix19_En18 
    input [18:0] Wgt_3_232, // sfix19_En18 
    input [18:0] Wgt_3_233, // sfix19_En18 
    input [18:0] Wgt_3_234, // sfix19_En18 
    input [18:0] Wgt_3_235, // sfix19_En18 
    input [18:0] Wgt_3_236, // sfix19_En18 
    input [18:0] Wgt_3_237, // sfix19_En18 
    input [18:0] Wgt_3_238, // sfix19_En18 
    input [18:0] Wgt_3_239, // sfix19_En18 
    input [18:0] Wgt_3_240, // sfix19_En18 
    input [18:0] Wgt_3_241, // sfix19_En18 
    input [18:0] Wgt_3_242, // sfix19_En18 
    input [18:0] Wgt_3_243, // sfix19_En18 
    input [18:0] Wgt_3_244, // sfix19_En18 
    input [18:0] Wgt_3_245, // sfix19_En18 
    input [18:0] Wgt_3_246, // sfix19_En18 
    input [18:0] Wgt_3_247, // sfix19_En18 
    input [18:0] Wgt_3_248, // sfix19_En18 
    input [18:0] Wgt_3_249, // sfix19_En18 
    input [18:0] Wgt_3_250, // sfix19_En18 
    input [18:0] Wgt_3_251, // sfix19_En18 
    input [18:0] Wgt_3_252, // sfix19_En18 
    input [18:0] Wgt_3_253, // sfix19_En18 
    input [18:0] Wgt_3_254, // sfix19_En18 
    input [18:0] Wgt_3_255, // sfix19_En18 
    input [18:0] Wgt_3_256, // sfix19_En18 
    input [18:0] Wgt_3_257, // sfix19_En18 
    input [18:0] Wgt_3_258, // sfix19_En18 
    input [18:0] Wgt_3_259, // sfix19_En18 
    input [18:0] Wgt_3_260, // sfix19_En18 
    input [18:0] Wgt_3_261, // sfix19_En18 
    input [18:0] Wgt_3_262, // sfix19_En18 
    input [18:0] Wgt_3_263, // sfix19_En18 
    input [18:0] Wgt_3_264, // sfix19_En18 
    input [18:0] Wgt_3_265, // sfix19_En18 
    input [18:0] Wgt_3_266, // sfix19_En18 
    input [18:0] Wgt_3_267, // sfix19_En18 
    input [18:0] Wgt_3_268, // sfix19_En18 
    input [18:0] Wgt_3_269, // sfix19_En18 
    input [18:0] Wgt_3_270, // sfix19_En18 
    input [18:0] Wgt_3_271, // sfix19_En18 
    input [18:0] Wgt_3_272, // sfix19_En18 
    input [18:0] Wgt_3_273, // sfix19_En18 
    input [18:0] Wgt_3_274, // sfix19_En18 
    input [18:0] Wgt_3_275, // sfix19_En18 
    input [18:0] Wgt_3_276, // sfix19_En18 
    input [18:0] Wgt_3_277, // sfix19_En18 
    input [18:0] Wgt_3_278, // sfix19_En18 
    input [18:0] Wgt_3_279, // sfix19_En18 
    input [18:0] Wgt_3_280, // sfix19_En18 
    input [18:0] Wgt_3_281, // sfix19_En18 
    input [18:0] Wgt_3_282, // sfix19_En18 
    input [18:0] Wgt_3_283, // sfix19_En18 
    input [18:0] Wgt_3_284, // sfix19_En18 
    input [18:0] Wgt_3_285, // sfix19_En18 
    input [18:0] Wgt_3_286, // sfix19_En18 
    input [18:0] Wgt_3_287, // sfix19_En18 
    input [18:0] Wgt_3_288, // sfix19_En18 
    input [18:0] Wgt_3_289, // sfix19_En18 
    input [18:0] Wgt_3_290, // sfix19_En18 
    input [18:0] Wgt_3_291, // sfix19_En18 
    input [18:0] Wgt_3_292, // sfix19_En18 
    input [18:0] Wgt_3_293, // sfix19_En18 
    input [18:0] Wgt_3_294, // sfix19_En18 
    input [18:0] Wgt_3_295, // sfix19_En18 
    input [18:0] Wgt_3_296, // sfix19_En18 
    input [18:0] Wgt_3_297, // sfix19_En18 
    input [18:0] Wgt_3_298, // sfix19_En18 
    input [18:0] Wgt_3_299, // sfix19_En18 
    input [18:0] Wgt_3_300, // sfix19_En18 
    input [18:0] Wgt_3_301, // sfix19_En18 
    input [18:0] Wgt_3_302, // sfix19_En18 
    input [18:0] Wgt_3_303, // sfix19_En18 
    input [18:0] Wgt_3_304, // sfix19_En18 
    input [18:0] Wgt_3_305, // sfix19_En18 
    input [18:0] Wgt_3_306, // sfix19_En18 
    input [18:0] Wgt_3_307, // sfix19_En18 
    input [18:0] Wgt_3_308, // sfix19_En18 
    input [18:0] Wgt_3_309, // sfix19_En18 
    input [18:0] Wgt_3_310, // sfix19_En18 
    input [18:0] Wgt_3_311, // sfix19_En18 
    input [18:0] Wgt_3_312, // sfix19_En18 
    input [18:0] Wgt_3_313, // sfix19_En18 
    input [18:0] Wgt_3_314, // sfix19_En18 
    input [18:0] Wgt_3_315, // sfix19_En18 
    input [18:0] Wgt_3_316, // sfix19_En18 
    input [18:0] Wgt_3_317, // sfix19_En18 
    input [18:0] Wgt_3_318, // sfix19_En18 
    input [18:0] Wgt_3_319, // sfix19_En18 
    input [18:0] Wgt_3_320, // sfix19_En18 
    input [18:0] Wgt_3_321, // sfix19_En18 
    input [18:0] Wgt_3_322, // sfix19_En18 
    input [18:0] Wgt_3_323, // sfix19_En18 
    input [18:0] Wgt_3_324, // sfix19_En18 
    input [18:0] Wgt_3_325, // sfix19_En18 
    input [18:0] Wgt_3_326, // sfix19_En18 
    input [18:0] Wgt_3_327, // sfix19_En18 
    input [18:0] Wgt_3_328, // sfix19_En18 
    input [18:0] Wgt_3_329, // sfix19_En18 
    input [18:0] Wgt_3_330, // sfix19_En18 
    input [18:0] Wgt_3_331, // sfix19_En18 
    input [18:0] Wgt_3_332, // sfix19_En18 
    input [18:0] Wgt_3_333, // sfix19_En18 
    input [18:0] Wgt_3_334, // sfix19_En18 
    input [18:0] Wgt_3_335, // sfix19_En18 
    input [18:0] Wgt_3_336, // sfix19_En18 
    input [18:0] Wgt_3_337, // sfix19_En18 
    input [18:0] Wgt_3_338, // sfix19_En18 
    input [18:0] Wgt_3_339, // sfix19_En18 
    input [18:0] Wgt_3_340, // sfix19_En18 
    input [18:0] Wgt_3_341, // sfix19_En18 
    input [18:0] Wgt_3_342, // sfix19_En18 
    input [18:0] Wgt_3_343, // sfix19_En18 
    input [18:0] Wgt_3_344, // sfix19_En18 
    input [18:0] Wgt_3_345, // sfix19_En18 
    input [18:0] Wgt_3_346, // sfix19_En18 
    input [18:0] Wgt_3_347, // sfix19_En18 
    input [18:0] Wgt_3_348, // sfix19_En18 
    input [18:0] Wgt_3_349, // sfix19_En18 
    input [18:0] Wgt_3_350, // sfix19_En18 
    input [18:0] Wgt_3_351, // sfix19_En18 
    input [18:0] Wgt_3_352, // sfix19_En18 
    input [18:0] Wgt_3_353, // sfix19_En18 
    input [18:0] Wgt_3_354, // sfix19_En18 
    input [18:0] Wgt_3_355, // sfix19_En18 
    input [18:0] Wgt_3_356, // sfix19_En18 
    input [18:0] Wgt_3_357, // sfix19_En18 
    input [18:0] Wgt_3_358, // sfix19_En18 
    input [18:0] Wgt_3_359, // sfix19_En18 
    input [18:0] Wgt_3_360, // sfix19_En18 
    input [18:0] Wgt_3_361, // sfix19_En18 
    input [18:0] Wgt_3_362, // sfix19_En18 
    input [18:0] Wgt_3_363, // sfix19_En18 
    input [18:0] Wgt_3_364, // sfix19_En18 
    input [18:0] Wgt_3_365, // sfix19_En18 
    input [18:0] Wgt_3_366, // sfix19_En18 
    input [18:0] Wgt_3_367, // sfix19_En18 
    input [18:0] Wgt_3_368, // sfix19_En18 
    input [18:0] Wgt_3_369, // sfix19_En18 
    input [18:0] Wgt_3_370, // sfix19_En18 
    input [18:0] Wgt_3_371, // sfix19_En18 
    input [18:0] Wgt_3_372, // sfix19_En18 
    input [18:0] Wgt_3_373, // sfix19_En18 
    input [18:0] Wgt_3_374, // sfix19_En18 
    input [18:0] Wgt_3_375, // sfix19_En18 
    input [18:0] Wgt_3_376, // sfix19_En18 
    input [18:0] Wgt_3_377, // sfix19_En18 
    input [18:0] Wgt_3_378, // sfix19_En18 
    input [18:0] Wgt_3_379, // sfix19_En18 
    input [18:0] Wgt_3_380, // sfix19_En18 
    input [18:0] Wgt_3_381, // sfix19_En18 
    input [18:0] Wgt_3_382, // sfix19_En18 
    input [18:0] Wgt_3_383, // sfix19_En18 
    input [18:0] Wgt_3_384, // sfix19_En18 
    input [18:0] Wgt_3_385, // sfix19_En18 
    input [18:0] Wgt_3_386, // sfix19_En18 
    input [18:0] Wgt_3_387, // sfix19_En18 
    input [18:0] Wgt_3_388, // sfix19_En18 
    input [18:0] Wgt_3_389, // sfix19_En18 
    input [18:0] Wgt_3_390, // sfix19_En18 
    input [18:0] Wgt_3_391, // sfix19_En18 
    input [18:0] Wgt_3_392, // sfix19_En18 
    input [18:0] Wgt_3_393, // sfix19_En18 
    input [18:0] Wgt_3_394, // sfix19_En18 
    input [18:0] Wgt_3_395, // sfix19_En18 
    input [18:0] Wgt_3_396, // sfix19_En18 
    input [18:0] Wgt_3_397, // sfix19_En18 
    input [18:0] Wgt_3_398, // sfix19_En18 
    input [18:0] Wgt_3_399, // sfix19_En18 
    input [18:0] Wgt_3_400, // sfix19_En18 
    input [18:0] Wgt_3_401, // sfix19_En18 
    input [18:0] Wgt_3_402, // sfix19_En18 
    input [18:0] Wgt_3_403, // sfix19_En18 
    input [18:0] Wgt_3_404, // sfix19_En18 
    input [18:0] Wgt_3_405, // sfix19_En18 
    input [18:0] Wgt_3_406, // sfix19_En18 
    input [18:0] Wgt_3_407, // sfix19_En18 
    input [18:0] Wgt_3_408, // sfix19_En18 
    input [18:0] Wgt_3_409, // sfix19_En18 
    input [18:0] Wgt_3_410, // sfix19_En18 
    input [18:0] Wgt_3_411, // sfix19_En18 
    input [18:0] Wgt_3_412, // sfix19_En18 
    input [18:0] Wgt_3_413, // sfix19_En18 
    input [18:0] Wgt_3_414, // sfix19_En18 
    input [18:0] Wgt_3_415, // sfix19_En18 
    input [18:0] Wgt_3_416, // sfix19_En18 
    input [18:0] Wgt_3_417, // sfix19_En18 
    input [18:0] Wgt_3_418, // sfix19_En18 
    input [18:0] Wgt_3_419, // sfix19_En18 
    input [18:0] Wgt_3_420, // sfix19_En18 
    input [18:0] Wgt_3_421, // sfix19_En18 
    input [18:0] Wgt_3_422, // sfix19_En18 
    input [18:0] Wgt_3_423, // sfix19_En18 
    input [18:0] Wgt_3_424, // sfix19_En18 
    input [18:0] Wgt_3_425, // sfix19_En18 
    input [18:0] Wgt_3_426, // sfix19_En18 
    input [18:0] Wgt_3_427, // sfix19_En18 
    input [18:0] Wgt_3_428, // sfix19_En18 
    input [18:0] Wgt_3_429, // sfix19_En18 
    input [18:0] Wgt_3_430, // sfix19_En18 
    input [18:0] Wgt_3_431, // sfix19_En18 
    input [18:0] Wgt_3_432, // sfix19_En18 
    input [18:0] Wgt_3_433, // sfix19_En18 
    input [18:0] Wgt_3_434, // sfix19_En18 
    input [18:0] Wgt_3_435, // sfix19_En18 
    input [18:0] Wgt_3_436, // sfix19_En18 
    input [18:0] Wgt_3_437, // sfix19_En18 
    input [18:0] Wgt_3_438, // sfix19_En18 
    input [18:0] Wgt_3_439, // sfix19_En18 
    input [18:0] Wgt_3_440, // sfix19_En18 
    input [18:0] Wgt_3_441, // sfix19_En18 
    input [18:0] Wgt_3_442, // sfix19_En18 
    input [18:0] Wgt_3_443, // sfix19_En18 
    input [18:0] Wgt_3_444, // sfix19_En18 
    input [18:0] Wgt_3_445, // sfix19_En18 
    input [18:0] Wgt_3_446, // sfix19_En18 
    input [18:0] Wgt_3_447, // sfix19_En18 
    input [18:0] Wgt_3_448, // sfix19_En18 
    input [18:0] Wgt_3_449, // sfix19_En18 
    input [18:0] Wgt_3_450, // sfix19_En18 
    input [18:0] Wgt_3_451, // sfix19_En18 
    input [18:0] Wgt_3_452, // sfix19_En18 
    input [18:0] Wgt_3_453, // sfix19_En18 
    input [18:0] Wgt_3_454, // sfix19_En18 
    input [18:0] Wgt_3_455, // sfix19_En18 
    input [18:0] Wgt_3_456, // sfix19_En18 
    input [18:0] Wgt_3_457, // sfix19_En18 
    input [18:0] Wgt_3_458, // sfix19_En18 
    input [18:0] Wgt_3_459, // sfix19_En18 
    input [18:0] Wgt_3_460, // sfix19_En18 
    input [18:0] Wgt_3_461, // sfix19_En18 
    input [18:0] Wgt_3_462, // sfix19_En18 
    input [18:0] Wgt_3_463, // sfix19_En18 
    input [18:0] Wgt_3_464, // sfix19_En18 
    input [18:0] Wgt_3_465, // sfix19_En18 
    input [18:0] Wgt_3_466, // sfix19_En18 
    input [18:0] Wgt_3_467, // sfix19_En18 
    input [18:0] Wgt_3_468, // sfix19_En18 
    input [18:0] Wgt_3_469, // sfix19_En18 
    input [18:0] Wgt_3_470, // sfix19_En18 
    input [18:0] Wgt_3_471, // sfix19_En18 
    input [18:0] Wgt_3_472, // sfix19_En18 
    input [18:0] Wgt_3_473, // sfix19_En18 
    input [18:0] Wgt_3_474, // sfix19_En18 
    input [18:0] Wgt_3_475, // sfix19_En18 
    input [18:0] Wgt_3_476, // sfix19_En18 
    input [18:0] Wgt_3_477, // sfix19_En18 
    input [18:0] Wgt_3_478, // sfix19_En18 
    input [18:0] Wgt_3_479, // sfix19_En18 
    input [18:0] Wgt_3_480, // sfix19_En18 
    input [18:0] Wgt_3_481, // sfix19_En18 
    input [18:0] Wgt_3_482, // sfix19_En18 
    input [18:0] Wgt_3_483, // sfix19_En18 
    input [18:0] Wgt_3_484, // sfix19_En18 
    input [18:0] Wgt_3_485, // sfix19_En18 
    input [18:0] Wgt_3_486, // sfix19_En18 
    input [18:0] Wgt_3_487, // sfix19_En18 
    input [18:0] Wgt_3_488, // sfix19_En18 
    input [18:0] Wgt_3_489, // sfix19_En18 
    input [18:0] Wgt_3_490, // sfix19_En18 
    input [18:0] Wgt_3_491, // sfix19_En18 
    input [18:0] Wgt_3_492, // sfix19_En18 
    input [18:0] Wgt_3_493, // sfix19_En18 
    input [18:0] Wgt_3_494, // sfix19_En18 
    input [18:0] Wgt_3_495, // sfix19_En18 
    input [18:0] Wgt_3_496, // sfix19_En18 
    input [18:0] Wgt_3_497, // sfix19_En18 
    input [18:0] Wgt_3_498, // sfix19_En18 
    input [18:0] Wgt_3_499, // sfix19_En18 
    input [18:0] Wgt_3_500, // sfix19_En18 
    input [18:0] Wgt_3_501, // sfix19_En18 
    input [18:0] Wgt_3_502, // sfix19_En18 
    input [18:0] Wgt_3_503, // sfix19_En18 
    input [18:0] Wgt_3_504, // sfix19_En18 
    input [18:0] Wgt_3_505, // sfix19_En18 
    input [18:0] Wgt_3_506, // sfix19_En18 
    input [18:0] Wgt_3_507, // sfix19_En18 
    input [18:0] Wgt_3_508, // sfix19_En18 
    input [18:0] Wgt_3_509, // sfix19_En18 
    input [18:0] Wgt_3_510, // sfix19_En18 
    input [18:0] Wgt_3_511, // sfix19_En18 
    input [18:0] Wgt_3_512, // sfix19_En18 
    input [18:0] Wgt_3_513, // sfix19_En18 
    input [18:0] Wgt_3_514, // sfix19_En18 
    input [18:0] Wgt_3_515, // sfix19_En18 
    input [18:0] Wgt_3_516, // sfix19_En18 
    input [18:0] Wgt_3_517, // sfix19_En18 
    input [18:0] Wgt_3_518, // sfix19_En18 
    input [18:0] Wgt_3_519, // sfix19_En18 
    input [18:0] Wgt_3_520, // sfix19_En18 
    input [18:0] Wgt_3_521, // sfix19_En18 
    input [18:0] Wgt_3_522, // sfix19_En18 
    input [18:0] Wgt_3_523, // sfix19_En18 
    input [18:0] Wgt_3_524, // sfix19_En18 
    input [18:0] Wgt_3_525, // sfix19_En18 
    input [18:0] Wgt_3_526, // sfix19_En18 
    input [18:0] Wgt_3_527, // sfix19_En18 
    input [18:0] Wgt_3_528, // sfix19_En18 
    input [18:0] Wgt_3_529, // sfix19_En18 
    input [18:0] Wgt_3_530, // sfix19_En18 
    input [18:0] Wgt_3_531, // sfix19_En18 
    input [18:0] Wgt_3_532, // sfix19_En18 
    input [18:0] Wgt_3_533, // sfix19_En18 
    input [18:0] Wgt_3_534, // sfix19_En18 
    input [18:0] Wgt_3_535, // sfix19_En18 
    input [18:0] Wgt_3_536, // sfix19_En18 
    input [18:0] Wgt_3_537, // sfix19_En18 
    input [18:0] Wgt_3_538, // sfix19_En18 
    input [18:0] Wgt_3_539, // sfix19_En18 
    input [18:0] Wgt_3_540, // sfix19_En18 
    input [18:0] Wgt_3_541, // sfix19_En18 
    input [18:0] Wgt_3_542, // sfix19_En18 
    input [18:0] Wgt_3_543, // sfix19_En18 
    input [18:0] Wgt_3_544, // sfix19_En18 
    input [18:0] Wgt_3_545, // sfix19_En18 
    input [18:0] Wgt_3_546, // sfix19_En18 
    input [18:0] Wgt_3_547, // sfix19_En18 
    input [18:0] Wgt_3_548, // sfix19_En18 
    input [18:0] Wgt_3_549, // sfix19_En18 
    input [18:0] Wgt_3_550, // sfix19_En18 
    input [18:0] Wgt_3_551, // sfix19_En18 
    input [18:0] Wgt_3_552, // sfix19_En18 
    input [18:0] Wgt_3_553, // sfix19_En18 
    input [18:0] Wgt_3_554, // sfix19_En18 
    input [18:0] Wgt_3_555, // sfix19_En18 
    input [18:0] Wgt_3_556, // sfix19_En18 
    input [18:0] Wgt_3_557, // sfix19_En18 
    input [18:0] Wgt_3_558, // sfix19_En18 
    input [18:0] Wgt_3_559, // sfix19_En18 
    input [18:0] Wgt_3_560, // sfix19_En18 
    input [18:0] Wgt_3_561, // sfix19_En18 
    input [18:0] Wgt_3_562, // sfix19_En18 
    input [18:0] Wgt_3_563, // sfix19_En18 
    input [18:0] Wgt_3_564, // sfix19_En18 
    input [18:0] Wgt_3_565, // sfix19_En18 
    input [18:0] Wgt_3_566, // sfix19_En18 
    input [18:0] Wgt_3_567, // sfix19_En18 
    input [18:0] Wgt_3_568, // sfix19_En18 
    input [18:0] Wgt_3_569, // sfix19_En18 
    input [18:0] Wgt_3_570, // sfix19_En18 
    input [18:0] Wgt_3_571, // sfix19_En18 
    input [18:0] Wgt_3_572, // sfix19_En18 
    input [18:0] Wgt_3_573, // sfix19_En18 
    input [18:0] Wgt_3_574, // sfix19_En18 
    input [18:0] Wgt_3_575, // sfix19_En18 
    input [18:0] Wgt_3_576, // sfix19_En18 
    input [18:0] Wgt_3_577, // sfix19_En18 
    input [18:0] Wgt_3_578, // sfix19_En18 
    input [18:0] Wgt_3_579, // sfix19_En18 
    input [18:0] Wgt_3_580, // sfix19_En18 
    input [18:0] Wgt_3_581, // sfix19_En18 
    input [18:0] Wgt_3_582, // sfix19_En18 
    input [18:0] Wgt_3_583, // sfix19_En18 
    input [18:0] Wgt_3_584, // sfix19_En18 
    input [18:0] Wgt_3_585, // sfix19_En18 
    input [18:0] Wgt_3_586, // sfix19_En18 
    input [18:0] Wgt_3_587, // sfix19_En18 
    input [18:0] Wgt_3_588, // sfix19_En18 
    input [18:0] Wgt_3_589, // sfix19_En18 
    input [18:0] Wgt_3_590, // sfix19_En18 
    input [18:0] Wgt_3_591, // sfix19_En18 
    input [18:0] Wgt_3_592, // sfix19_En18 
    input [18:0] Wgt_3_593, // sfix19_En18 
    input [18:0] Wgt_3_594, // sfix19_En18 
    input [18:0] Wgt_3_595, // sfix19_En18 
    input [18:0] Wgt_3_596, // sfix19_En18 
    input [18:0] Wgt_3_597, // sfix19_En18 
    input [18:0] Wgt_3_598, // sfix19_En18 
    input [18:0] Wgt_3_599, // sfix19_En18 
    input [18:0] Wgt_3_600, // sfix19_En18 
    input [18:0] Wgt_3_601, // sfix19_En18 
    input [18:0] Wgt_3_602, // sfix19_En18 
    input [18:0] Wgt_3_603, // sfix19_En18 
    input [18:0] Wgt_3_604, // sfix19_En18 
    input [18:0] Wgt_3_605, // sfix19_En18 
    input [18:0] Wgt_3_606, // sfix19_En18 
    input [18:0] Wgt_3_607, // sfix19_En18 
    input [18:0] Wgt_3_608, // sfix19_En18 
    input [18:0] Wgt_3_609, // sfix19_En18 
    input [18:0] Wgt_3_610, // sfix19_En18 
    input [18:0] Wgt_3_611, // sfix19_En18 
    input [18:0] Wgt_3_612, // sfix19_En18 
    input [18:0] Wgt_3_613, // sfix19_En18 
    input [18:0] Wgt_3_614, // sfix19_En18 
    input [18:0] Wgt_3_615, // sfix19_En18 
    input [18:0] Wgt_3_616, // sfix19_En18 
    input [18:0] Wgt_3_617, // sfix19_En18 
    input [18:0] Wgt_3_618, // sfix19_En18 
    input [18:0] Wgt_3_619, // sfix19_En18 
    input [18:0] Wgt_3_620, // sfix19_En18 
    input [18:0] Wgt_3_621, // sfix19_En18 
    input [18:0] Wgt_3_622, // sfix19_En18 
    input [18:0] Wgt_3_623, // sfix19_En18 
    input [18:0] Wgt_3_624, // sfix19_En18 
    input [18:0] Wgt_3_625, // sfix19_En18 
    input [18:0] Wgt_3_626, // sfix19_En18 
    input [18:0] Wgt_3_627, // sfix19_En18 
    input [18:0] Wgt_3_628, // sfix19_En18 
    input [18:0] Wgt_3_629, // sfix19_En18 
    input [18:0] Wgt_3_630, // sfix19_En18 
    input [18:0] Wgt_3_631, // sfix19_En18 
    input [18:0] Wgt_3_632, // sfix19_En18 
    input [18:0] Wgt_3_633, // sfix19_En18 
    input [18:0] Wgt_3_634, // sfix19_En18 
    input [18:0] Wgt_3_635, // sfix19_En18 
    input [18:0] Wgt_3_636, // sfix19_En18 
    input [18:0] Wgt_3_637, // sfix19_En18 
    input [18:0] Wgt_3_638, // sfix19_En18 
    input [18:0] Wgt_3_639, // sfix19_En18 
    input [18:0] Wgt_3_640, // sfix19_En18 
    input [18:0] Wgt_3_641, // sfix19_En18 
    input [18:0] Wgt_3_642, // sfix19_En18 
    input [18:0] Wgt_3_643, // sfix19_En18 
    input [18:0] Wgt_3_644, // sfix19_En18 
    input [18:0] Wgt_3_645, // sfix19_En18 
    input [18:0] Wgt_3_646, // sfix19_En18 
    input [18:0] Wgt_3_647, // sfix19_En18 
    input [18:0] Wgt_3_648, // sfix19_En18 
    input [18:0] Wgt_3_649, // sfix19_En18 
    input [18:0] Wgt_3_650, // sfix19_En18 
    input [18:0] Wgt_3_651, // sfix19_En18 
    input [18:0] Wgt_3_652, // sfix19_En18 
    input [18:0] Wgt_3_653, // sfix19_En18 
    input [18:0] Wgt_3_654, // sfix19_En18 
    input [18:0] Wgt_3_655, // sfix19_En18 
    input [18:0] Wgt_3_656, // sfix19_En18 
    input [18:0] Wgt_3_657, // sfix19_En18 
    input [18:0] Wgt_3_658, // sfix19_En18 
    input [18:0] Wgt_3_659, // sfix19_En18 
    input [18:0] Wgt_3_660, // sfix19_En18 
    input [18:0] Wgt_3_661, // sfix19_En18 
    input [18:0] Wgt_3_662, // sfix19_En18 
    input [18:0] Wgt_3_663, // sfix19_En18 
    input [18:0] Wgt_3_664, // sfix19_En18 
    input [18:0] Wgt_3_665, // sfix19_En18 
    input [18:0] Wgt_3_666, // sfix19_En18 
    input [18:0] Wgt_3_667, // sfix19_En18 
    input [18:0] Wgt_3_668, // sfix19_En18 
    input [18:0] Wgt_3_669, // sfix19_En18 
    input [18:0] Wgt_3_670, // sfix19_En18 
    input [18:0] Wgt_3_671, // sfix19_En18 
    input [18:0] Wgt_3_672, // sfix19_En18 
    input [18:0] Wgt_3_673, // sfix19_En18 
    input [18:0] Wgt_3_674, // sfix19_En18 
    input [18:0] Wgt_3_675, // sfix19_En18 
    input [18:0] Wgt_3_676, // sfix19_En18 
    input [18:0] Wgt_3_677, // sfix19_En18 
    input [18:0] Wgt_3_678, // sfix19_En18 
    input [18:0] Wgt_3_679, // sfix19_En18 
    input [18:0] Wgt_3_680, // sfix19_En18 
    input [18:0] Wgt_3_681, // sfix19_En18 
    input [18:0] Wgt_3_682, // sfix19_En18 
    input [18:0] Wgt_3_683, // sfix19_En18 
    input [18:0] Wgt_3_684, // sfix19_En18 
    input [18:0] Wgt_3_685, // sfix19_En18 
    input [18:0] Wgt_3_686, // sfix19_En18 
    input [18:0] Wgt_3_687, // sfix19_En18 
    input [18:0] Wgt_3_688, // sfix19_En18 
    input [18:0] Wgt_3_689, // sfix19_En18 
    input [18:0] Wgt_3_690, // sfix19_En18 
    input [18:0] Wgt_3_691, // sfix19_En18 
    input [18:0] Wgt_3_692, // sfix19_En18 
    input [18:0] Wgt_3_693, // sfix19_En18 
    input [18:0] Wgt_3_694, // sfix19_En18 
    input [18:0] Wgt_3_695, // sfix19_En18 
    input [18:0] Wgt_3_696, // sfix19_En18 
    input [18:0] Wgt_3_697, // sfix19_En18 
    input [18:0] Wgt_3_698, // sfix19_En18 
    input [18:0] Wgt_3_699, // sfix19_En18 
    input [18:0] Wgt_3_700, // sfix19_En18 
    input [18:0] Wgt_3_701, // sfix19_En18 
    input [18:0] Wgt_3_702, // sfix19_En18 
    input [18:0] Wgt_3_703, // sfix19_En18 
    input [18:0] Wgt_3_704, // sfix19_En18 
    input [18:0] Wgt_3_705, // sfix19_En18 
    input [18:0] Wgt_3_706, // sfix19_En18 
    input [18:0] Wgt_3_707, // sfix19_En18 
    input [18:0] Wgt_3_708, // sfix19_En18 
    input [18:0] Wgt_3_709, // sfix19_En18 
    input [18:0] Wgt_3_710, // sfix19_En18 
    input [18:0] Wgt_3_711, // sfix19_En18 
    input [18:0] Wgt_3_712, // sfix19_En18 
    input [18:0] Wgt_3_713, // sfix19_En18 
    input [18:0] Wgt_3_714, // sfix19_En18 
    input [18:0] Wgt_3_715, // sfix19_En18 
    input [18:0] Wgt_3_716, // sfix19_En18 
    input [18:0] Wgt_3_717, // sfix19_En18 
    input [18:0] Wgt_3_718, // sfix19_En18 
    input [18:0] Wgt_3_719, // sfix19_En18 
    input [18:0] Wgt_3_720, // sfix19_En18 
    input [18:0] Wgt_3_721, // sfix19_En18 
    input [18:0] Wgt_3_722, // sfix19_En18 
    input [18:0] Wgt_3_723, // sfix19_En18 
    input [18:0] Wgt_3_724, // sfix19_En18 
    input [18:0] Wgt_3_725, // sfix19_En18 
    input [18:0] Wgt_3_726, // sfix19_En18 
    input [18:0] Wgt_3_727, // sfix19_En18 
    input [18:0] Wgt_3_728, // sfix19_En18 
    input [18:0] Wgt_3_729, // sfix19_En18 
    input [18:0] Wgt_3_730, // sfix19_En18 
    input [18:0] Wgt_3_731, // sfix19_En18 
    input [18:0] Wgt_3_732, // sfix19_En18 
    input [18:0] Wgt_3_733, // sfix19_En18 
    input [18:0] Wgt_3_734, // sfix19_En18 
    input [18:0] Wgt_3_735, // sfix19_En18 
    input [18:0] Wgt_3_736, // sfix19_En18 
    input [18:0] Wgt_3_737, // sfix19_En18 
    input [18:0] Wgt_3_738, // sfix19_En18 
    input [18:0] Wgt_3_739, // sfix19_En18 
    input [18:0] Wgt_3_740, // sfix19_En18 
    input [18:0] Wgt_3_741, // sfix19_En18 
    input [18:0] Wgt_3_742, // sfix19_En18 
    input [18:0] Wgt_3_743, // sfix19_En18 
    input [18:0] Wgt_3_744, // sfix19_En18 
    input [18:0] Wgt_3_745, // sfix19_En18 
    input [18:0] Wgt_3_746, // sfix19_En18 
    input [18:0] Wgt_3_747, // sfix19_En18 
    input [18:0] Wgt_3_748, // sfix19_En18 
    input [18:0] Wgt_3_749, // sfix19_En18 
    input [18:0] Wgt_3_750, // sfix19_En18 
    input [18:0] Wgt_3_751, // sfix19_En18 
    input [18:0] Wgt_3_752, // sfix19_En18 
    input [18:0] Wgt_3_753, // sfix19_En18 
    input [18:0] Wgt_3_754, // sfix19_En18 
    input [18:0] Wgt_3_755, // sfix19_En18 
    input [18:0] Wgt_3_756, // sfix19_En18 
    input [18:0] Wgt_3_757, // sfix19_En18 
    input [18:0] Wgt_3_758, // sfix19_En18 
    input [18:0] Wgt_3_759, // sfix19_En18 
    input [18:0] Wgt_3_760, // sfix19_En18 
    input [18:0] Wgt_3_761, // sfix19_En18 
    input [18:0] Wgt_3_762, // sfix19_En18 
    input [18:0] Wgt_3_763, // sfix19_En18 
    input [18:0] Wgt_3_764, // sfix19_En18 
    input [18:0] Wgt_3_765, // sfix19_En18 
    input [18:0] Wgt_3_766, // sfix19_En18 
    input [18:0] Wgt_3_767, // sfix19_En18 
    input [18:0] Wgt_3_768, // sfix19_En18 
    input [18:0] Wgt_3_769, // sfix19_En18 
    input [18:0] Wgt_3_770, // sfix19_En18 
    input [18:0] Wgt_3_771, // sfix19_En18 
    input [18:0] Wgt_3_772, // sfix19_En18 
    input [18:0] Wgt_3_773, // sfix19_En18 
    input [18:0] Wgt_3_774, // sfix19_En18 
    input [18:0] Wgt_3_775, // sfix19_En18 
    input [18:0] Wgt_3_776, // sfix19_En18 
    input [18:0] Wgt_3_777, // sfix19_En18 
    input [18:0] Wgt_3_778, // sfix19_En18 
    input [18:0] Wgt_3_779, // sfix19_En18 
    input [18:0] Wgt_3_780, // sfix19_En18 
    input [18:0] Wgt_3_781, // sfix19_En18 
    input [18:0] Wgt_3_782, // sfix19_En18 
    input [18:0] Wgt_3_783, // sfix19_En18 
    input [18:0] Wgt_3_784, // sfix19_En18 
    input [18:0] Wgt_4_0, // sfix19_En18 
    input [18:0] Wgt_4_1, // sfix19_En18 
    input [18:0] Wgt_4_2, // sfix19_En18 
    input [18:0] Wgt_4_3, // sfix19_En18 
    input [18:0] Wgt_4_4, // sfix19_En18 
    input [18:0] Wgt_4_5, // sfix19_En18 
    input [18:0] Wgt_4_6, // sfix19_En18 
    input [18:0] Wgt_4_7, // sfix19_En18 
    input [18:0] Wgt_4_8, // sfix19_En18 
    input [18:0] Wgt_4_9, // sfix19_En18 
    input [18:0] Wgt_4_10, // sfix19_En18 
    input [18:0] Wgt_4_11, // sfix19_En18 
    input [18:0] Wgt_4_12, // sfix19_En18 
    input [18:0] Wgt_4_13, // sfix19_En18 
    input [18:0] Wgt_4_14, // sfix19_En18 
    input [18:0] Wgt_4_15, // sfix19_En18 
    input [18:0] Wgt_4_16, // sfix19_En18 
    input [18:0] Wgt_4_17, // sfix19_En18 
    input [18:0] Wgt_4_18, // sfix19_En18 
    input [18:0] Wgt_4_19, // sfix19_En18 
    input [18:0] Wgt_4_20, // sfix19_En18 
    input [18:0] Wgt_4_21, // sfix19_En18 
    input [18:0] Wgt_4_22, // sfix19_En18 
    input [18:0] Wgt_4_23, // sfix19_En18 
    input [18:0] Wgt_4_24, // sfix19_En18 
    input [18:0] Wgt_4_25, // sfix19_En18 
    input [18:0] Wgt_4_26, // sfix19_En18 
    input [18:0] Wgt_4_27, // sfix19_En18 
    input [18:0] Wgt_4_28, // sfix19_En18 
    input [18:0] Wgt_4_29, // sfix19_En18 
    input [18:0] Wgt_4_30, // sfix19_En18 
    input [18:0] Wgt_4_31, // sfix19_En18 
    input [18:0] Wgt_4_32, // sfix19_En18 
    input [18:0] Wgt_4_33, // sfix19_En18 
    input [18:0] Wgt_4_34, // sfix19_En18 
    input [18:0] Wgt_4_35, // sfix19_En18 
    input [18:0] Wgt_4_36, // sfix19_En18 
    input [18:0] Wgt_4_37, // sfix19_En18 
    input [18:0] Wgt_4_38, // sfix19_En18 
    input [18:0] Wgt_4_39, // sfix19_En18 
    input [18:0] Wgt_4_40, // sfix19_En18 
    input [18:0] Wgt_4_41, // sfix19_En18 
    input [18:0] Wgt_4_42, // sfix19_En18 
    input [18:0] Wgt_4_43, // sfix19_En18 
    input [18:0] Wgt_4_44, // sfix19_En18 
    input [18:0] Wgt_4_45, // sfix19_En18 
    input [18:0] Wgt_4_46, // sfix19_En18 
    input [18:0] Wgt_4_47, // sfix19_En18 
    input [18:0] Wgt_4_48, // sfix19_En18 
    input [18:0] Wgt_4_49, // sfix19_En18 
    input [18:0] Wgt_4_50, // sfix19_En18 
    input [18:0] Wgt_4_51, // sfix19_En18 
    input [18:0] Wgt_4_52, // sfix19_En18 
    input [18:0] Wgt_4_53, // sfix19_En18 
    input [18:0] Wgt_4_54, // sfix19_En18 
    input [18:0] Wgt_4_55, // sfix19_En18 
    input [18:0] Wgt_4_56, // sfix19_En18 
    input [18:0] Wgt_4_57, // sfix19_En18 
    input [18:0] Wgt_4_58, // sfix19_En18 
    input [18:0] Wgt_4_59, // sfix19_En18 
    input [18:0] Wgt_4_60, // sfix19_En18 
    input [18:0] Wgt_4_61, // sfix19_En18 
    input [18:0] Wgt_4_62, // sfix19_En18 
    input [18:0] Wgt_4_63, // sfix19_En18 
    input [18:0] Wgt_4_64, // sfix19_En18 
    input [18:0] Wgt_4_65, // sfix19_En18 
    input [18:0] Wgt_4_66, // sfix19_En18 
    input [18:0] Wgt_4_67, // sfix19_En18 
    input [18:0] Wgt_4_68, // sfix19_En18 
    input [18:0] Wgt_4_69, // sfix19_En18 
    input [18:0] Wgt_4_70, // sfix19_En18 
    input [18:0] Wgt_4_71, // sfix19_En18 
    input [18:0] Wgt_4_72, // sfix19_En18 
    input [18:0] Wgt_4_73, // sfix19_En18 
    input [18:0] Wgt_4_74, // sfix19_En18 
    input [18:0] Wgt_4_75, // sfix19_En18 
    input [18:0] Wgt_4_76, // sfix19_En18 
    input [18:0] Wgt_4_77, // sfix19_En18 
    input [18:0] Wgt_4_78, // sfix19_En18 
    input [18:0] Wgt_4_79, // sfix19_En18 
    input [18:0] Wgt_4_80, // sfix19_En18 
    input [18:0] Wgt_4_81, // sfix19_En18 
    input [18:0] Wgt_4_82, // sfix19_En18 
    input [18:0] Wgt_4_83, // sfix19_En18 
    input [18:0] Wgt_4_84, // sfix19_En18 
    input [18:0] Wgt_4_85, // sfix19_En18 
    input [18:0] Wgt_4_86, // sfix19_En18 
    input [18:0] Wgt_4_87, // sfix19_En18 
    input [18:0] Wgt_4_88, // sfix19_En18 
    input [18:0] Wgt_4_89, // sfix19_En18 
    input [18:0] Wgt_4_90, // sfix19_En18 
    input [18:0] Wgt_4_91, // sfix19_En18 
    input [18:0] Wgt_4_92, // sfix19_En18 
    input [18:0] Wgt_4_93, // sfix19_En18 
    input [18:0] Wgt_4_94, // sfix19_En18 
    input [18:0] Wgt_4_95, // sfix19_En18 
    input [18:0] Wgt_4_96, // sfix19_En18 
    input [18:0] Wgt_4_97, // sfix19_En18 
    input [18:0] Wgt_4_98, // sfix19_En18 
    input [18:0] Wgt_4_99, // sfix19_En18 
    input [18:0] Wgt_4_100, // sfix19_En18 
    input [18:0] Wgt_4_101, // sfix19_En18 
    input [18:0] Wgt_4_102, // sfix19_En18 
    input [18:0] Wgt_4_103, // sfix19_En18 
    input [18:0] Wgt_4_104, // sfix19_En18 
    input [18:0] Wgt_4_105, // sfix19_En18 
    input [18:0] Wgt_4_106, // sfix19_En18 
    input [18:0] Wgt_4_107, // sfix19_En18 
    input [18:0] Wgt_4_108, // sfix19_En18 
    input [18:0] Wgt_4_109, // sfix19_En18 
    input [18:0] Wgt_4_110, // sfix19_En18 
    input [18:0] Wgt_4_111, // sfix19_En18 
    input [18:0] Wgt_4_112, // sfix19_En18 
    input [18:0] Wgt_4_113, // sfix19_En18 
    input [18:0] Wgt_4_114, // sfix19_En18 
    input [18:0] Wgt_4_115, // sfix19_En18 
    input [18:0] Wgt_4_116, // sfix19_En18 
    input [18:0] Wgt_4_117, // sfix19_En18 
    input [18:0] Wgt_4_118, // sfix19_En18 
    input [18:0] Wgt_4_119, // sfix19_En18 
    input [18:0] Wgt_4_120, // sfix19_En18 
    input [18:0] Wgt_4_121, // sfix19_En18 
    input [18:0] Wgt_4_122, // sfix19_En18 
    input [18:0] Wgt_4_123, // sfix19_En18 
    input [18:0] Wgt_4_124, // sfix19_En18 
    input [18:0] Wgt_4_125, // sfix19_En18 
    input [18:0] Wgt_4_126, // sfix19_En18 
    input [18:0] Wgt_4_127, // sfix19_En18 
    input [18:0] Wgt_4_128, // sfix19_En18 
    input [18:0] Wgt_4_129, // sfix19_En18 
    input [18:0] Wgt_4_130, // sfix19_En18 
    input [18:0] Wgt_4_131, // sfix19_En18 
    input [18:0] Wgt_4_132, // sfix19_En18 
    input [18:0] Wgt_4_133, // sfix19_En18 
    input [18:0] Wgt_4_134, // sfix19_En18 
    input [18:0] Wgt_4_135, // sfix19_En18 
    input [18:0] Wgt_4_136, // sfix19_En18 
    input [18:0] Wgt_4_137, // sfix19_En18 
    input [18:0] Wgt_4_138, // sfix19_En18 
    input [18:0] Wgt_4_139, // sfix19_En18 
    input [18:0] Wgt_4_140, // sfix19_En18 
    input [18:0] Wgt_4_141, // sfix19_En18 
    input [18:0] Wgt_4_142, // sfix19_En18 
    input [18:0] Wgt_4_143, // sfix19_En18 
    input [18:0] Wgt_4_144, // sfix19_En18 
    input [18:0] Wgt_4_145, // sfix19_En18 
    input [18:0] Wgt_4_146, // sfix19_En18 
    input [18:0] Wgt_4_147, // sfix19_En18 
    input [18:0] Wgt_4_148, // sfix19_En18 
    input [18:0] Wgt_4_149, // sfix19_En18 
    input [18:0] Wgt_4_150, // sfix19_En18 
    input [18:0] Wgt_4_151, // sfix19_En18 
    input [18:0] Wgt_4_152, // sfix19_En18 
    input [18:0] Wgt_4_153, // sfix19_En18 
    input [18:0] Wgt_4_154, // sfix19_En18 
    input [18:0] Wgt_4_155, // sfix19_En18 
    input [18:0] Wgt_4_156, // sfix19_En18 
    input [18:0] Wgt_4_157, // sfix19_En18 
    input [18:0] Wgt_4_158, // sfix19_En18 
    input [18:0] Wgt_4_159, // sfix19_En18 
    input [18:0] Wgt_4_160, // sfix19_En18 
    input [18:0] Wgt_4_161, // sfix19_En18 
    input [18:0] Wgt_4_162, // sfix19_En18 
    input [18:0] Wgt_4_163, // sfix19_En18 
    input [18:0] Wgt_4_164, // sfix19_En18 
    input [18:0] Wgt_4_165, // sfix19_En18 
    input [18:0] Wgt_4_166, // sfix19_En18 
    input [18:0] Wgt_4_167, // sfix19_En18 
    input [18:0] Wgt_4_168, // sfix19_En18 
    input [18:0] Wgt_4_169, // sfix19_En18 
    input [18:0] Wgt_4_170, // sfix19_En18 
    input [18:0] Wgt_4_171, // sfix19_En18 
    input [18:0] Wgt_4_172, // sfix19_En18 
    input [18:0] Wgt_4_173, // sfix19_En18 
    input [18:0] Wgt_4_174, // sfix19_En18 
    input [18:0] Wgt_4_175, // sfix19_En18 
    input [18:0] Wgt_4_176, // sfix19_En18 
    input [18:0] Wgt_4_177, // sfix19_En18 
    input [18:0] Wgt_4_178, // sfix19_En18 
    input [18:0] Wgt_4_179, // sfix19_En18 
    input [18:0] Wgt_4_180, // sfix19_En18 
    input [18:0] Wgt_4_181, // sfix19_En18 
    input [18:0] Wgt_4_182, // sfix19_En18 
    input [18:0] Wgt_4_183, // sfix19_En18 
    input [18:0] Wgt_4_184, // sfix19_En18 
    input [18:0] Wgt_4_185, // sfix19_En18 
    input [18:0] Wgt_4_186, // sfix19_En18 
    input [18:0] Wgt_4_187, // sfix19_En18 
    input [18:0] Wgt_4_188, // sfix19_En18 
    input [18:0] Wgt_4_189, // sfix19_En18 
    input [18:0] Wgt_4_190, // sfix19_En18 
    input [18:0] Wgt_4_191, // sfix19_En18 
    input [18:0] Wgt_4_192, // sfix19_En18 
    input [18:0] Wgt_4_193, // sfix19_En18 
    input [18:0] Wgt_4_194, // sfix19_En18 
    input [18:0] Wgt_4_195, // sfix19_En18 
    input [18:0] Wgt_4_196, // sfix19_En18 
    input [18:0] Wgt_4_197, // sfix19_En18 
    input [18:0] Wgt_4_198, // sfix19_En18 
    input [18:0] Wgt_4_199, // sfix19_En18 
    input [18:0] Wgt_4_200, // sfix19_En18 
    input [18:0] Wgt_4_201, // sfix19_En18 
    input [18:0] Wgt_4_202, // sfix19_En18 
    input [18:0] Wgt_4_203, // sfix19_En18 
    input [18:0] Wgt_4_204, // sfix19_En18 
    input [18:0] Wgt_4_205, // sfix19_En18 
    input [18:0] Wgt_4_206, // sfix19_En18 
    input [18:0] Wgt_4_207, // sfix19_En18 
    input [18:0] Wgt_4_208, // sfix19_En18 
    input [18:0] Wgt_4_209, // sfix19_En18 
    input [18:0] Wgt_4_210, // sfix19_En18 
    input [18:0] Wgt_4_211, // sfix19_En18 
    input [18:0] Wgt_4_212, // sfix19_En18 
    input [18:0] Wgt_4_213, // sfix19_En18 
    input [18:0] Wgt_4_214, // sfix19_En18 
    input [18:0] Wgt_4_215, // sfix19_En18 
    input [18:0] Wgt_4_216, // sfix19_En18 
    input [18:0] Wgt_4_217, // sfix19_En18 
    input [18:0] Wgt_4_218, // sfix19_En18 
    input [18:0] Wgt_4_219, // sfix19_En18 
    input [18:0] Wgt_4_220, // sfix19_En18 
    input [18:0] Wgt_4_221, // sfix19_En18 
    input [18:0] Wgt_4_222, // sfix19_En18 
    input [18:0] Wgt_4_223, // sfix19_En18 
    input [18:0] Wgt_4_224, // sfix19_En18 
    input [18:0] Wgt_4_225, // sfix19_En18 
    input [18:0] Wgt_4_226, // sfix19_En18 
    input [18:0] Wgt_4_227, // sfix19_En18 
    input [18:0] Wgt_4_228, // sfix19_En18 
    input [18:0] Wgt_4_229, // sfix19_En18 
    input [18:0] Wgt_4_230, // sfix19_En18 
    input [18:0] Wgt_4_231, // sfix19_En18 
    input [18:0] Wgt_4_232, // sfix19_En18 
    input [18:0] Wgt_4_233, // sfix19_En18 
    input [18:0] Wgt_4_234, // sfix19_En18 
    input [18:0] Wgt_4_235, // sfix19_En18 
    input [18:0] Wgt_4_236, // sfix19_En18 
    input [18:0] Wgt_4_237, // sfix19_En18 
    input [18:0] Wgt_4_238, // sfix19_En18 
    input [18:0] Wgt_4_239, // sfix19_En18 
    input [18:0] Wgt_4_240, // sfix19_En18 
    input [18:0] Wgt_4_241, // sfix19_En18 
    input [18:0] Wgt_4_242, // sfix19_En18 
    input [18:0] Wgt_4_243, // sfix19_En18 
    input [18:0] Wgt_4_244, // sfix19_En18 
    input [18:0] Wgt_4_245, // sfix19_En18 
    input [18:0] Wgt_4_246, // sfix19_En18 
    input [18:0] Wgt_4_247, // sfix19_En18 
    input [18:0] Wgt_4_248, // sfix19_En18 
    input [18:0] Wgt_4_249, // sfix19_En18 
    input [18:0] Wgt_4_250, // sfix19_En18 
    input [18:0] Wgt_4_251, // sfix19_En18 
    input [18:0] Wgt_4_252, // sfix19_En18 
    input [18:0] Wgt_4_253, // sfix19_En18 
    input [18:0] Wgt_4_254, // sfix19_En18 
    input [18:0] Wgt_4_255, // sfix19_En18 
    input [18:0] Wgt_4_256, // sfix19_En18 
    input [18:0] Wgt_4_257, // sfix19_En18 
    input [18:0] Wgt_4_258, // sfix19_En18 
    input [18:0] Wgt_4_259, // sfix19_En18 
    input [18:0] Wgt_4_260, // sfix19_En18 
    input [18:0] Wgt_4_261, // sfix19_En18 
    input [18:0] Wgt_4_262, // sfix19_En18 
    input [18:0] Wgt_4_263, // sfix19_En18 
    input [18:0] Wgt_4_264, // sfix19_En18 
    input [18:0] Wgt_4_265, // sfix19_En18 
    input [18:0] Wgt_4_266, // sfix19_En18 
    input [18:0] Wgt_4_267, // sfix19_En18 
    input [18:0] Wgt_4_268, // sfix19_En18 
    input [18:0] Wgt_4_269, // sfix19_En18 
    input [18:0] Wgt_4_270, // sfix19_En18 
    input [18:0] Wgt_4_271, // sfix19_En18 
    input [18:0] Wgt_4_272, // sfix19_En18 
    input [18:0] Wgt_4_273, // sfix19_En18 
    input [18:0] Wgt_4_274, // sfix19_En18 
    input [18:0] Wgt_4_275, // sfix19_En18 
    input [18:0] Wgt_4_276, // sfix19_En18 
    input [18:0] Wgt_4_277, // sfix19_En18 
    input [18:0] Wgt_4_278, // sfix19_En18 
    input [18:0] Wgt_4_279, // sfix19_En18 
    input [18:0] Wgt_4_280, // sfix19_En18 
    input [18:0] Wgt_4_281, // sfix19_En18 
    input [18:0] Wgt_4_282, // sfix19_En18 
    input [18:0] Wgt_4_283, // sfix19_En18 
    input [18:0] Wgt_4_284, // sfix19_En18 
    input [18:0] Wgt_4_285, // sfix19_En18 
    input [18:0] Wgt_4_286, // sfix19_En18 
    input [18:0] Wgt_4_287, // sfix19_En18 
    input [18:0] Wgt_4_288, // sfix19_En18 
    input [18:0] Wgt_4_289, // sfix19_En18 
    input [18:0] Wgt_4_290, // sfix19_En18 
    input [18:0] Wgt_4_291, // sfix19_En18 
    input [18:0] Wgt_4_292, // sfix19_En18 
    input [18:0] Wgt_4_293, // sfix19_En18 
    input [18:0] Wgt_4_294, // sfix19_En18 
    input [18:0] Wgt_4_295, // sfix19_En18 
    input [18:0] Wgt_4_296, // sfix19_En18 
    input [18:0] Wgt_4_297, // sfix19_En18 
    input [18:0] Wgt_4_298, // sfix19_En18 
    input [18:0] Wgt_4_299, // sfix19_En18 
    input [18:0] Wgt_4_300, // sfix19_En18 
    input [18:0] Wgt_4_301, // sfix19_En18 
    input [18:0] Wgt_4_302, // sfix19_En18 
    input [18:0] Wgt_4_303, // sfix19_En18 
    input [18:0] Wgt_4_304, // sfix19_En18 
    input [18:0] Wgt_4_305, // sfix19_En18 
    input [18:0] Wgt_4_306, // sfix19_En18 
    input [18:0] Wgt_4_307, // sfix19_En18 
    input [18:0] Wgt_4_308, // sfix19_En18 
    input [18:0] Wgt_4_309, // sfix19_En18 
    input [18:0] Wgt_4_310, // sfix19_En18 
    input [18:0] Wgt_4_311, // sfix19_En18 
    input [18:0] Wgt_4_312, // sfix19_En18 
    input [18:0] Wgt_4_313, // sfix19_En18 
    input [18:0] Wgt_4_314, // sfix19_En18 
    input [18:0] Wgt_4_315, // sfix19_En18 
    input [18:0] Wgt_4_316, // sfix19_En18 
    input [18:0] Wgt_4_317, // sfix19_En18 
    input [18:0] Wgt_4_318, // sfix19_En18 
    input [18:0] Wgt_4_319, // sfix19_En18 
    input [18:0] Wgt_4_320, // sfix19_En18 
    input [18:0] Wgt_4_321, // sfix19_En18 
    input [18:0] Wgt_4_322, // sfix19_En18 
    input [18:0] Wgt_4_323, // sfix19_En18 
    input [18:0] Wgt_4_324, // sfix19_En18 
    input [18:0] Wgt_4_325, // sfix19_En18 
    input [18:0] Wgt_4_326, // sfix19_En18 
    input [18:0] Wgt_4_327, // sfix19_En18 
    input [18:0] Wgt_4_328, // sfix19_En18 
    input [18:0] Wgt_4_329, // sfix19_En18 
    input [18:0] Wgt_4_330, // sfix19_En18 
    input [18:0] Wgt_4_331, // sfix19_En18 
    input [18:0] Wgt_4_332, // sfix19_En18 
    input [18:0] Wgt_4_333, // sfix19_En18 
    input [18:0] Wgt_4_334, // sfix19_En18 
    input [18:0] Wgt_4_335, // sfix19_En18 
    input [18:0] Wgt_4_336, // sfix19_En18 
    input [18:0] Wgt_4_337, // sfix19_En18 
    input [18:0] Wgt_4_338, // sfix19_En18 
    input [18:0] Wgt_4_339, // sfix19_En18 
    input [18:0] Wgt_4_340, // sfix19_En18 
    input [18:0] Wgt_4_341, // sfix19_En18 
    input [18:0] Wgt_4_342, // sfix19_En18 
    input [18:0] Wgt_4_343, // sfix19_En18 
    input [18:0] Wgt_4_344, // sfix19_En18 
    input [18:0] Wgt_4_345, // sfix19_En18 
    input [18:0] Wgt_4_346, // sfix19_En18 
    input [18:0] Wgt_4_347, // sfix19_En18 
    input [18:0] Wgt_4_348, // sfix19_En18 
    input [18:0] Wgt_4_349, // sfix19_En18 
    input [18:0] Wgt_4_350, // sfix19_En18 
    input [18:0] Wgt_4_351, // sfix19_En18 
    input [18:0] Wgt_4_352, // sfix19_En18 
    input [18:0] Wgt_4_353, // sfix19_En18 
    input [18:0] Wgt_4_354, // sfix19_En18 
    input [18:0] Wgt_4_355, // sfix19_En18 
    input [18:0] Wgt_4_356, // sfix19_En18 
    input [18:0] Wgt_4_357, // sfix19_En18 
    input [18:0] Wgt_4_358, // sfix19_En18 
    input [18:0] Wgt_4_359, // sfix19_En18 
    input [18:0] Wgt_4_360, // sfix19_En18 
    input [18:0] Wgt_4_361, // sfix19_En18 
    input [18:0] Wgt_4_362, // sfix19_En18 
    input [18:0] Wgt_4_363, // sfix19_En18 
    input [18:0] Wgt_4_364, // sfix19_En18 
    input [18:0] Wgt_4_365, // sfix19_En18 
    input [18:0] Wgt_4_366, // sfix19_En18 
    input [18:0] Wgt_4_367, // sfix19_En18 
    input [18:0] Wgt_4_368, // sfix19_En18 
    input [18:0] Wgt_4_369, // sfix19_En18 
    input [18:0] Wgt_4_370, // sfix19_En18 
    input [18:0] Wgt_4_371, // sfix19_En18 
    input [18:0] Wgt_4_372, // sfix19_En18 
    input [18:0] Wgt_4_373, // sfix19_En18 
    input [18:0] Wgt_4_374, // sfix19_En18 
    input [18:0] Wgt_4_375, // sfix19_En18 
    input [18:0] Wgt_4_376, // sfix19_En18 
    input [18:0] Wgt_4_377, // sfix19_En18 
    input [18:0] Wgt_4_378, // sfix19_En18 
    input [18:0] Wgt_4_379, // sfix19_En18 
    input [18:0] Wgt_4_380, // sfix19_En18 
    input [18:0] Wgt_4_381, // sfix19_En18 
    input [18:0] Wgt_4_382, // sfix19_En18 
    input [18:0] Wgt_4_383, // sfix19_En18 
    input [18:0] Wgt_4_384, // sfix19_En18 
    input [18:0] Wgt_4_385, // sfix19_En18 
    input [18:0] Wgt_4_386, // sfix19_En18 
    input [18:0] Wgt_4_387, // sfix19_En18 
    input [18:0] Wgt_4_388, // sfix19_En18 
    input [18:0] Wgt_4_389, // sfix19_En18 
    input [18:0] Wgt_4_390, // sfix19_En18 
    input [18:0] Wgt_4_391, // sfix19_En18 
    input [18:0] Wgt_4_392, // sfix19_En18 
    input [18:0] Wgt_4_393, // sfix19_En18 
    input [18:0] Wgt_4_394, // sfix19_En18 
    input [18:0] Wgt_4_395, // sfix19_En18 
    input [18:0] Wgt_4_396, // sfix19_En18 
    input [18:0] Wgt_4_397, // sfix19_En18 
    input [18:0] Wgt_4_398, // sfix19_En18 
    input [18:0] Wgt_4_399, // sfix19_En18 
    input [18:0] Wgt_4_400, // sfix19_En18 
    input [18:0] Wgt_4_401, // sfix19_En18 
    input [18:0] Wgt_4_402, // sfix19_En18 
    input [18:0] Wgt_4_403, // sfix19_En18 
    input [18:0] Wgt_4_404, // sfix19_En18 
    input [18:0] Wgt_4_405, // sfix19_En18 
    input [18:0] Wgt_4_406, // sfix19_En18 
    input [18:0] Wgt_4_407, // sfix19_En18 
    input [18:0] Wgt_4_408, // sfix19_En18 
    input [18:0] Wgt_4_409, // sfix19_En18 
    input [18:0] Wgt_4_410, // sfix19_En18 
    input [18:0] Wgt_4_411, // sfix19_En18 
    input [18:0] Wgt_4_412, // sfix19_En18 
    input [18:0] Wgt_4_413, // sfix19_En18 
    input [18:0] Wgt_4_414, // sfix19_En18 
    input [18:0] Wgt_4_415, // sfix19_En18 
    input [18:0] Wgt_4_416, // sfix19_En18 
    input [18:0] Wgt_4_417, // sfix19_En18 
    input [18:0] Wgt_4_418, // sfix19_En18 
    input [18:0] Wgt_4_419, // sfix19_En18 
    input [18:0] Wgt_4_420, // sfix19_En18 
    input [18:0] Wgt_4_421, // sfix19_En18 
    input [18:0] Wgt_4_422, // sfix19_En18 
    input [18:0] Wgt_4_423, // sfix19_En18 
    input [18:0] Wgt_4_424, // sfix19_En18 
    input [18:0] Wgt_4_425, // sfix19_En18 
    input [18:0] Wgt_4_426, // sfix19_En18 
    input [18:0] Wgt_4_427, // sfix19_En18 
    input [18:0] Wgt_4_428, // sfix19_En18 
    input [18:0] Wgt_4_429, // sfix19_En18 
    input [18:0] Wgt_4_430, // sfix19_En18 
    input [18:0] Wgt_4_431, // sfix19_En18 
    input [18:0] Wgt_4_432, // sfix19_En18 
    input [18:0] Wgt_4_433, // sfix19_En18 
    input [18:0] Wgt_4_434, // sfix19_En18 
    input [18:0] Wgt_4_435, // sfix19_En18 
    input [18:0] Wgt_4_436, // sfix19_En18 
    input [18:0] Wgt_4_437, // sfix19_En18 
    input [18:0] Wgt_4_438, // sfix19_En18 
    input [18:0] Wgt_4_439, // sfix19_En18 
    input [18:0] Wgt_4_440, // sfix19_En18 
    input [18:0] Wgt_4_441, // sfix19_En18 
    input [18:0] Wgt_4_442, // sfix19_En18 
    input [18:0] Wgt_4_443, // sfix19_En18 
    input [18:0] Wgt_4_444, // sfix19_En18 
    input [18:0] Wgt_4_445, // sfix19_En18 
    input [18:0] Wgt_4_446, // sfix19_En18 
    input [18:0] Wgt_4_447, // sfix19_En18 
    input [18:0] Wgt_4_448, // sfix19_En18 
    input [18:0] Wgt_4_449, // sfix19_En18 
    input [18:0] Wgt_4_450, // sfix19_En18 
    input [18:0] Wgt_4_451, // sfix19_En18 
    input [18:0] Wgt_4_452, // sfix19_En18 
    input [18:0] Wgt_4_453, // sfix19_En18 
    input [18:0] Wgt_4_454, // sfix19_En18 
    input [18:0] Wgt_4_455, // sfix19_En18 
    input [18:0] Wgt_4_456, // sfix19_En18 
    input [18:0] Wgt_4_457, // sfix19_En18 
    input [18:0] Wgt_4_458, // sfix19_En18 
    input [18:0] Wgt_4_459, // sfix19_En18 
    input [18:0] Wgt_4_460, // sfix19_En18 
    input [18:0] Wgt_4_461, // sfix19_En18 
    input [18:0] Wgt_4_462, // sfix19_En18 
    input [18:0] Wgt_4_463, // sfix19_En18 
    input [18:0] Wgt_4_464, // sfix19_En18 
    input [18:0] Wgt_4_465, // sfix19_En18 
    input [18:0] Wgt_4_466, // sfix19_En18 
    input [18:0] Wgt_4_467, // sfix19_En18 
    input [18:0] Wgt_4_468, // sfix19_En18 
    input [18:0] Wgt_4_469, // sfix19_En18 
    input [18:0] Wgt_4_470, // sfix19_En18 
    input [18:0] Wgt_4_471, // sfix19_En18 
    input [18:0] Wgt_4_472, // sfix19_En18 
    input [18:0] Wgt_4_473, // sfix19_En18 
    input [18:0] Wgt_4_474, // sfix19_En18 
    input [18:0] Wgt_4_475, // sfix19_En18 
    input [18:0] Wgt_4_476, // sfix19_En18 
    input [18:0] Wgt_4_477, // sfix19_En18 
    input [18:0] Wgt_4_478, // sfix19_En18 
    input [18:0] Wgt_4_479, // sfix19_En18 
    input [18:0] Wgt_4_480, // sfix19_En18 
    input [18:0] Wgt_4_481, // sfix19_En18 
    input [18:0] Wgt_4_482, // sfix19_En18 
    input [18:0] Wgt_4_483, // sfix19_En18 
    input [18:0] Wgt_4_484, // sfix19_En18 
    input [18:0] Wgt_4_485, // sfix19_En18 
    input [18:0] Wgt_4_486, // sfix19_En18 
    input [18:0] Wgt_4_487, // sfix19_En18 
    input [18:0] Wgt_4_488, // sfix19_En18 
    input [18:0] Wgt_4_489, // sfix19_En18 
    input [18:0] Wgt_4_490, // sfix19_En18 
    input [18:0] Wgt_4_491, // sfix19_En18 
    input [18:0] Wgt_4_492, // sfix19_En18 
    input [18:0] Wgt_4_493, // sfix19_En18 
    input [18:0] Wgt_4_494, // sfix19_En18 
    input [18:0] Wgt_4_495, // sfix19_En18 
    input [18:0] Wgt_4_496, // sfix19_En18 
    input [18:0] Wgt_4_497, // sfix19_En18 
    input [18:0] Wgt_4_498, // sfix19_En18 
    input [18:0] Wgt_4_499, // sfix19_En18 
    input [18:0] Wgt_4_500, // sfix19_En18 
    input [18:0] Wgt_4_501, // sfix19_En18 
    input [18:0] Wgt_4_502, // sfix19_En18 
    input [18:0] Wgt_4_503, // sfix19_En18 
    input [18:0] Wgt_4_504, // sfix19_En18 
    input [18:0] Wgt_4_505, // sfix19_En18 
    input [18:0] Wgt_4_506, // sfix19_En18 
    input [18:0] Wgt_4_507, // sfix19_En18 
    input [18:0] Wgt_4_508, // sfix19_En18 
    input [18:0] Wgt_4_509, // sfix19_En18 
    input [18:0] Wgt_4_510, // sfix19_En18 
    input [18:0] Wgt_4_511, // sfix19_En18 
    input [18:0] Wgt_4_512, // sfix19_En18 
    input [18:0] Wgt_4_513, // sfix19_En18 
    input [18:0] Wgt_4_514, // sfix19_En18 
    input [18:0] Wgt_4_515, // sfix19_En18 
    input [18:0] Wgt_4_516, // sfix19_En18 
    input [18:0] Wgt_4_517, // sfix19_En18 
    input [18:0] Wgt_4_518, // sfix19_En18 
    input [18:0] Wgt_4_519, // sfix19_En18 
    input [18:0] Wgt_4_520, // sfix19_En18 
    input [18:0] Wgt_4_521, // sfix19_En18 
    input [18:0] Wgt_4_522, // sfix19_En18 
    input [18:0] Wgt_4_523, // sfix19_En18 
    input [18:0] Wgt_4_524, // sfix19_En18 
    input [18:0] Wgt_4_525, // sfix19_En18 
    input [18:0] Wgt_4_526, // sfix19_En18 
    input [18:0] Wgt_4_527, // sfix19_En18 
    input [18:0] Wgt_4_528, // sfix19_En18 
    input [18:0] Wgt_4_529, // sfix19_En18 
    input [18:0] Wgt_4_530, // sfix19_En18 
    input [18:0] Wgt_4_531, // sfix19_En18 
    input [18:0] Wgt_4_532, // sfix19_En18 
    input [18:0] Wgt_4_533, // sfix19_En18 
    input [18:0] Wgt_4_534, // sfix19_En18 
    input [18:0] Wgt_4_535, // sfix19_En18 
    input [18:0] Wgt_4_536, // sfix19_En18 
    input [18:0] Wgt_4_537, // sfix19_En18 
    input [18:0] Wgt_4_538, // sfix19_En18 
    input [18:0] Wgt_4_539, // sfix19_En18 
    input [18:0] Wgt_4_540, // sfix19_En18 
    input [18:0] Wgt_4_541, // sfix19_En18 
    input [18:0] Wgt_4_542, // sfix19_En18 
    input [18:0] Wgt_4_543, // sfix19_En18 
    input [18:0] Wgt_4_544, // sfix19_En18 
    input [18:0] Wgt_4_545, // sfix19_En18 
    input [18:0] Wgt_4_546, // sfix19_En18 
    input [18:0] Wgt_4_547, // sfix19_En18 
    input [18:0] Wgt_4_548, // sfix19_En18 
    input [18:0] Wgt_4_549, // sfix19_En18 
    input [18:0] Wgt_4_550, // sfix19_En18 
    input [18:0] Wgt_4_551, // sfix19_En18 
    input [18:0] Wgt_4_552, // sfix19_En18 
    input [18:0] Wgt_4_553, // sfix19_En18 
    input [18:0] Wgt_4_554, // sfix19_En18 
    input [18:0] Wgt_4_555, // sfix19_En18 
    input [18:0] Wgt_4_556, // sfix19_En18 
    input [18:0] Wgt_4_557, // sfix19_En18 
    input [18:0] Wgt_4_558, // sfix19_En18 
    input [18:0] Wgt_4_559, // sfix19_En18 
    input [18:0] Wgt_4_560, // sfix19_En18 
    input [18:0] Wgt_4_561, // sfix19_En18 
    input [18:0] Wgt_4_562, // sfix19_En18 
    input [18:0] Wgt_4_563, // sfix19_En18 
    input [18:0] Wgt_4_564, // sfix19_En18 
    input [18:0] Wgt_4_565, // sfix19_En18 
    input [18:0] Wgt_4_566, // sfix19_En18 
    input [18:0] Wgt_4_567, // sfix19_En18 
    input [18:0] Wgt_4_568, // sfix19_En18 
    input [18:0] Wgt_4_569, // sfix19_En18 
    input [18:0] Wgt_4_570, // sfix19_En18 
    input [18:0] Wgt_4_571, // sfix19_En18 
    input [18:0] Wgt_4_572, // sfix19_En18 
    input [18:0] Wgt_4_573, // sfix19_En18 
    input [18:0] Wgt_4_574, // sfix19_En18 
    input [18:0] Wgt_4_575, // sfix19_En18 
    input [18:0] Wgt_4_576, // sfix19_En18 
    input [18:0] Wgt_4_577, // sfix19_En18 
    input [18:0] Wgt_4_578, // sfix19_En18 
    input [18:0] Wgt_4_579, // sfix19_En18 
    input [18:0] Wgt_4_580, // sfix19_En18 
    input [18:0] Wgt_4_581, // sfix19_En18 
    input [18:0] Wgt_4_582, // sfix19_En18 
    input [18:0] Wgt_4_583, // sfix19_En18 
    input [18:0] Wgt_4_584, // sfix19_En18 
    input [18:0] Wgt_4_585, // sfix19_En18 
    input [18:0] Wgt_4_586, // sfix19_En18 
    input [18:0] Wgt_4_587, // sfix19_En18 
    input [18:0] Wgt_4_588, // sfix19_En18 
    input [18:0] Wgt_4_589, // sfix19_En18 
    input [18:0] Wgt_4_590, // sfix19_En18 
    input [18:0] Wgt_4_591, // sfix19_En18 
    input [18:0] Wgt_4_592, // sfix19_En18 
    input [18:0] Wgt_4_593, // sfix19_En18 
    input [18:0] Wgt_4_594, // sfix19_En18 
    input [18:0] Wgt_4_595, // sfix19_En18 
    input [18:0] Wgt_4_596, // sfix19_En18 
    input [18:0] Wgt_4_597, // sfix19_En18 
    input [18:0] Wgt_4_598, // sfix19_En18 
    input [18:0] Wgt_4_599, // sfix19_En18 
    input [18:0] Wgt_4_600, // sfix19_En18 
    input [18:0] Wgt_4_601, // sfix19_En18 
    input [18:0] Wgt_4_602, // sfix19_En18 
    input [18:0] Wgt_4_603, // sfix19_En18 
    input [18:0] Wgt_4_604, // sfix19_En18 
    input [18:0] Wgt_4_605, // sfix19_En18 
    input [18:0] Wgt_4_606, // sfix19_En18 
    input [18:0] Wgt_4_607, // sfix19_En18 
    input [18:0] Wgt_4_608, // sfix19_En18 
    input [18:0] Wgt_4_609, // sfix19_En18 
    input [18:0] Wgt_4_610, // sfix19_En18 
    input [18:0] Wgt_4_611, // sfix19_En18 
    input [18:0] Wgt_4_612, // sfix19_En18 
    input [18:0] Wgt_4_613, // sfix19_En18 
    input [18:0] Wgt_4_614, // sfix19_En18 
    input [18:0] Wgt_4_615, // sfix19_En18 
    input [18:0] Wgt_4_616, // sfix19_En18 
    input [18:0] Wgt_4_617, // sfix19_En18 
    input [18:0] Wgt_4_618, // sfix19_En18 
    input [18:0] Wgt_4_619, // sfix19_En18 
    input [18:0] Wgt_4_620, // sfix19_En18 
    input [18:0] Wgt_4_621, // sfix19_En18 
    input [18:0] Wgt_4_622, // sfix19_En18 
    input [18:0] Wgt_4_623, // sfix19_En18 
    input [18:0] Wgt_4_624, // sfix19_En18 
    input [18:0] Wgt_4_625, // sfix19_En18 
    input [18:0] Wgt_4_626, // sfix19_En18 
    input [18:0] Wgt_4_627, // sfix19_En18 
    input [18:0] Wgt_4_628, // sfix19_En18 
    input [18:0] Wgt_4_629, // sfix19_En18 
    input [18:0] Wgt_4_630, // sfix19_En18 
    input [18:0] Wgt_4_631, // sfix19_En18 
    input [18:0] Wgt_4_632, // sfix19_En18 
    input [18:0] Wgt_4_633, // sfix19_En18 
    input [18:0] Wgt_4_634, // sfix19_En18 
    input [18:0] Wgt_4_635, // sfix19_En18 
    input [18:0] Wgt_4_636, // sfix19_En18 
    input [18:0] Wgt_4_637, // sfix19_En18 
    input [18:0] Wgt_4_638, // sfix19_En18 
    input [18:0] Wgt_4_639, // sfix19_En18 
    input [18:0] Wgt_4_640, // sfix19_En18 
    input [18:0] Wgt_4_641, // sfix19_En18 
    input [18:0] Wgt_4_642, // sfix19_En18 
    input [18:0] Wgt_4_643, // sfix19_En18 
    input [18:0] Wgt_4_644, // sfix19_En18 
    input [18:0] Wgt_4_645, // sfix19_En18 
    input [18:0] Wgt_4_646, // sfix19_En18 
    input [18:0] Wgt_4_647, // sfix19_En18 
    input [18:0] Wgt_4_648, // sfix19_En18 
    input [18:0] Wgt_4_649, // sfix19_En18 
    input [18:0] Wgt_4_650, // sfix19_En18 
    input [18:0] Wgt_4_651, // sfix19_En18 
    input [18:0] Wgt_4_652, // sfix19_En18 
    input [18:0] Wgt_4_653, // sfix19_En18 
    input [18:0] Wgt_4_654, // sfix19_En18 
    input [18:0] Wgt_4_655, // sfix19_En18 
    input [18:0] Wgt_4_656, // sfix19_En18 
    input [18:0] Wgt_4_657, // sfix19_En18 
    input [18:0] Wgt_4_658, // sfix19_En18 
    input [18:0] Wgt_4_659, // sfix19_En18 
    input [18:0] Wgt_4_660, // sfix19_En18 
    input [18:0] Wgt_4_661, // sfix19_En18 
    input [18:0] Wgt_4_662, // sfix19_En18 
    input [18:0] Wgt_4_663, // sfix19_En18 
    input [18:0] Wgt_4_664, // sfix19_En18 
    input [18:0] Wgt_4_665, // sfix19_En18 
    input [18:0] Wgt_4_666, // sfix19_En18 
    input [18:0] Wgt_4_667, // sfix19_En18 
    input [18:0] Wgt_4_668, // sfix19_En18 
    input [18:0] Wgt_4_669, // sfix19_En18 
    input [18:0] Wgt_4_670, // sfix19_En18 
    input [18:0] Wgt_4_671, // sfix19_En18 
    input [18:0] Wgt_4_672, // sfix19_En18 
    input [18:0] Wgt_4_673, // sfix19_En18 
    input [18:0] Wgt_4_674, // sfix19_En18 
    input [18:0] Wgt_4_675, // sfix19_En18 
    input [18:0] Wgt_4_676, // sfix19_En18 
    input [18:0] Wgt_4_677, // sfix19_En18 
    input [18:0] Wgt_4_678, // sfix19_En18 
    input [18:0] Wgt_4_679, // sfix19_En18 
    input [18:0] Wgt_4_680, // sfix19_En18 
    input [18:0] Wgt_4_681, // sfix19_En18 
    input [18:0] Wgt_4_682, // sfix19_En18 
    input [18:0] Wgt_4_683, // sfix19_En18 
    input [18:0] Wgt_4_684, // sfix19_En18 
    input [18:0] Wgt_4_685, // sfix19_En18 
    input [18:0] Wgt_4_686, // sfix19_En18 
    input [18:0] Wgt_4_687, // sfix19_En18 
    input [18:0] Wgt_4_688, // sfix19_En18 
    input [18:0] Wgt_4_689, // sfix19_En18 
    input [18:0] Wgt_4_690, // sfix19_En18 
    input [18:0] Wgt_4_691, // sfix19_En18 
    input [18:0] Wgt_4_692, // sfix19_En18 
    input [18:0] Wgt_4_693, // sfix19_En18 
    input [18:0] Wgt_4_694, // sfix19_En18 
    input [18:0] Wgt_4_695, // sfix19_En18 
    input [18:0] Wgt_4_696, // sfix19_En18 
    input [18:0] Wgt_4_697, // sfix19_En18 
    input [18:0] Wgt_4_698, // sfix19_En18 
    input [18:0] Wgt_4_699, // sfix19_En18 
    input [18:0] Wgt_4_700, // sfix19_En18 
    input [18:0] Wgt_4_701, // sfix19_En18 
    input [18:0] Wgt_4_702, // sfix19_En18 
    input [18:0] Wgt_4_703, // sfix19_En18 
    input [18:0] Wgt_4_704, // sfix19_En18 
    input [18:0] Wgt_4_705, // sfix19_En18 
    input [18:0] Wgt_4_706, // sfix19_En18 
    input [18:0] Wgt_4_707, // sfix19_En18 
    input [18:0] Wgt_4_708, // sfix19_En18 
    input [18:0] Wgt_4_709, // sfix19_En18 
    input [18:0] Wgt_4_710, // sfix19_En18 
    input [18:0] Wgt_4_711, // sfix19_En18 
    input [18:0] Wgt_4_712, // sfix19_En18 
    input [18:0] Wgt_4_713, // sfix19_En18 
    input [18:0] Wgt_4_714, // sfix19_En18 
    input [18:0] Wgt_4_715, // sfix19_En18 
    input [18:0] Wgt_4_716, // sfix19_En18 
    input [18:0] Wgt_4_717, // sfix19_En18 
    input [18:0] Wgt_4_718, // sfix19_En18 
    input [18:0] Wgt_4_719, // sfix19_En18 
    input [18:0] Wgt_4_720, // sfix19_En18 
    input [18:0] Wgt_4_721, // sfix19_En18 
    input [18:0] Wgt_4_722, // sfix19_En18 
    input [18:0] Wgt_4_723, // sfix19_En18 
    input [18:0] Wgt_4_724, // sfix19_En18 
    input [18:0] Wgt_4_725, // sfix19_En18 
    input [18:0] Wgt_4_726, // sfix19_En18 
    input [18:0] Wgt_4_727, // sfix19_En18 
    input [18:0] Wgt_4_728, // sfix19_En18 
    input [18:0] Wgt_4_729, // sfix19_En18 
    input [18:0] Wgt_4_730, // sfix19_En18 
    input [18:0] Wgt_4_731, // sfix19_En18 
    input [18:0] Wgt_4_732, // sfix19_En18 
    input [18:0] Wgt_4_733, // sfix19_En18 
    input [18:0] Wgt_4_734, // sfix19_En18 
    input [18:0] Wgt_4_735, // sfix19_En18 
    input [18:0] Wgt_4_736, // sfix19_En18 
    input [18:0] Wgt_4_737, // sfix19_En18 
    input [18:0] Wgt_4_738, // sfix19_En18 
    input [18:0] Wgt_4_739, // sfix19_En18 
    input [18:0] Wgt_4_740, // sfix19_En18 
    input [18:0] Wgt_4_741, // sfix19_En18 
    input [18:0] Wgt_4_742, // sfix19_En18 
    input [18:0] Wgt_4_743, // sfix19_En18 
    input [18:0] Wgt_4_744, // sfix19_En18 
    input [18:0] Wgt_4_745, // sfix19_En18 
    input [18:0] Wgt_4_746, // sfix19_En18 
    input [18:0] Wgt_4_747, // sfix19_En18 
    input [18:0] Wgt_4_748, // sfix19_En18 
    input [18:0] Wgt_4_749, // sfix19_En18 
    input [18:0] Wgt_4_750, // sfix19_En18 
    input [18:0] Wgt_4_751, // sfix19_En18 
    input [18:0] Wgt_4_752, // sfix19_En18 
    input [18:0] Wgt_4_753, // sfix19_En18 
    input [18:0] Wgt_4_754, // sfix19_En18 
    input [18:0] Wgt_4_755, // sfix19_En18 
    input [18:0] Wgt_4_756, // sfix19_En18 
    input [18:0] Wgt_4_757, // sfix19_En18 
    input [18:0] Wgt_4_758, // sfix19_En18 
    input [18:0] Wgt_4_759, // sfix19_En18 
    input [18:0] Wgt_4_760, // sfix19_En18 
    input [18:0] Wgt_4_761, // sfix19_En18 
    input [18:0] Wgt_4_762, // sfix19_En18 
    input [18:0] Wgt_4_763, // sfix19_En18 
    input [18:0] Wgt_4_764, // sfix19_En18 
    input [18:0] Wgt_4_765, // sfix19_En18 
    input [18:0] Wgt_4_766, // sfix19_En18 
    input [18:0] Wgt_4_767, // sfix19_En18 
    input [18:0] Wgt_4_768, // sfix19_En18 
    input [18:0] Wgt_4_769, // sfix19_En18 
    input [18:0] Wgt_4_770, // sfix19_En18 
    input [18:0] Wgt_4_771, // sfix19_En18 
    input [18:0] Wgt_4_772, // sfix19_En18 
    input [18:0] Wgt_4_773, // sfix19_En18 
    input [18:0] Wgt_4_774, // sfix19_En18 
    input [18:0] Wgt_4_775, // sfix19_En18 
    input [18:0] Wgt_4_776, // sfix19_En18 
    input [18:0] Wgt_4_777, // sfix19_En18 
    input [18:0] Wgt_4_778, // sfix19_En18 
    input [18:0] Wgt_4_779, // sfix19_En18 
    input [18:0] Wgt_4_780, // sfix19_En18 
    input [18:0] Wgt_4_781, // sfix19_En18 
    input [18:0] Wgt_4_782, // sfix19_En18 
    input [18:0] Wgt_4_783, // sfix19_En18 
    input [18:0] Wgt_4_784, // sfix19_En18 
    input [18:0] Wgt_5_0, // sfix19_En18 
    input [18:0] Wgt_5_1, // sfix19_En18 
    input [18:0] Wgt_5_2, // sfix19_En18 
    input [18:0] Wgt_5_3, // sfix19_En18 
    input [18:0] Wgt_5_4, // sfix19_En18 
    input [18:0] Wgt_5_5, // sfix19_En18 
    input [18:0] Wgt_5_6, // sfix19_En18 
    input [18:0] Wgt_5_7, // sfix19_En18 
    input [18:0] Wgt_5_8, // sfix19_En18 
    input [18:0] Wgt_5_9, // sfix19_En18 
    input [18:0] Wgt_5_10, // sfix19_En18 
    input [18:0] Wgt_5_11, // sfix19_En18 
    input [18:0] Wgt_5_12, // sfix19_En18 
    input [18:0] Wgt_5_13, // sfix19_En18 
    input [18:0] Wgt_5_14, // sfix19_En18 
    input [18:0] Wgt_5_15, // sfix19_En18 
    input [18:0] Wgt_5_16, // sfix19_En18 
    input [18:0] Wgt_5_17, // sfix19_En18 
    input [18:0] Wgt_5_18, // sfix19_En18 
    input [18:0] Wgt_5_19, // sfix19_En18 
    input [18:0] Wgt_5_20, // sfix19_En18 
    input [18:0] Wgt_5_21, // sfix19_En18 
    input [18:0] Wgt_5_22, // sfix19_En18 
    input [18:0] Wgt_5_23, // sfix19_En18 
    input [18:0] Wgt_5_24, // sfix19_En18 
    input [18:0] Wgt_5_25, // sfix19_En18 
    input [18:0] Wgt_5_26, // sfix19_En18 
    input [18:0] Wgt_5_27, // sfix19_En18 
    input [18:0] Wgt_5_28, // sfix19_En18 
    input [18:0] Wgt_5_29, // sfix19_En18 
    input [18:0] Wgt_5_30, // sfix19_En18 
    input [18:0] Wgt_5_31, // sfix19_En18 
    input [18:0] Wgt_5_32, // sfix19_En18 
    input [18:0] Wgt_5_33, // sfix19_En18 
    input [18:0] Wgt_5_34, // sfix19_En18 
    input [18:0] Wgt_5_35, // sfix19_En18 
    input [18:0] Wgt_5_36, // sfix19_En18 
    input [18:0] Wgt_5_37, // sfix19_En18 
    input [18:0] Wgt_5_38, // sfix19_En18 
    input [18:0] Wgt_5_39, // sfix19_En18 
    input [18:0] Wgt_5_40, // sfix19_En18 
    input [18:0] Wgt_5_41, // sfix19_En18 
    input [18:0] Wgt_5_42, // sfix19_En18 
    input [18:0] Wgt_5_43, // sfix19_En18 
    input [18:0] Wgt_5_44, // sfix19_En18 
    input [18:0] Wgt_5_45, // sfix19_En18 
    input [18:0] Wgt_5_46, // sfix19_En18 
    input [18:0] Wgt_5_47, // sfix19_En18 
    input [18:0] Wgt_5_48, // sfix19_En18 
    input [18:0] Wgt_5_49, // sfix19_En18 
    input [18:0] Wgt_5_50, // sfix19_En18 
    input [18:0] Wgt_5_51, // sfix19_En18 
    input [18:0] Wgt_5_52, // sfix19_En18 
    input [18:0] Wgt_5_53, // sfix19_En18 
    input [18:0] Wgt_5_54, // sfix19_En18 
    input [18:0] Wgt_5_55, // sfix19_En18 
    input [18:0] Wgt_5_56, // sfix19_En18 
    input [18:0] Wgt_5_57, // sfix19_En18 
    input [18:0] Wgt_5_58, // sfix19_En18 
    input [18:0] Wgt_5_59, // sfix19_En18 
    input [18:0] Wgt_5_60, // sfix19_En18 
    input [18:0] Wgt_5_61, // sfix19_En18 
    input [18:0] Wgt_5_62, // sfix19_En18 
    input [18:0] Wgt_5_63, // sfix19_En18 
    input [18:0] Wgt_5_64, // sfix19_En18 
    input [18:0] Wgt_5_65, // sfix19_En18 
    input [18:0] Wgt_5_66, // sfix19_En18 
    input [18:0] Wgt_5_67, // sfix19_En18 
    input [18:0] Wgt_5_68, // sfix19_En18 
    input [18:0] Wgt_5_69, // sfix19_En18 
    input [18:0] Wgt_5_70, // sfix19_En18 
    input [18:0] Wgt_5_71, // sfix19_En18 
    input [18:0] Wgt_5_72, // sfix19_En18 
    input [18:0] Wgt_5_73, // sfix19_En18 
    input [18:0] Wgt_5_74, // sfix19_En18 
    input [18:0] Wgt_5_75, // sfix19_En18 
    input [18:0] Wgt_5_76, // sfix19_En18 
    input [18:0] Wgt_5_77, // sfix19_En18 
    input [18:0] Wgt_5_78, // sfix19_En18 
    input [18:0] Wgt_5_79, // sfix19_En18 
    input [18:0] Wgt_5_80, // sfix19_En18 
    input [18:0] Wgt_5_81, // sfix19_En18 
    input [18:0] Wgt_5_82, // sfix19_En18 
    input [18:0] Wgt_5_83, // sfix19_En18 
    input [18:0] Wgt_5_84, // sfix19_En18 
    input [18:0] Wgt_5_85, // sfix19_En18 
    input [18:0] Wgt_5_86, // sfix19_En18 
    input [18:0] Wgt_5_87, // sfix19_En18 
    input [18:0] Wgt_5_88, // sfix19_En18 
    input [18:0] Wgt_5_89, // sfix19_En18 
    input [18:0] Wgt_5_90, // sfix19_En18 
    input [18:0] Wgt_5_91, // sfix19_En18 
    input [18:0] Wgt_5_92, // sfix19_En18 
    input [18:0] Wgt_5_93, // sfix19_En18 
    input [18:0] Wgt_5_94, // sfix19_En18 
    input [18:0] Wgt_5_95, // sfix19_En18 
    input [18:0] Wgt_5_96, // sfix19_En18 
    input [18:0] Wgt_5_97, // sfix19_En18 
    input [18:0] Wgt_5_98, // sfix19_En18 
    input [18:0] Wgt_5_99, // sfix19_En18 
    input [18:0] Wgt_5_100, // sfix19_En18 
    input [18:0] Wgt_5_101, // sfix19_En18 
    input [18:0] Wgt_5_102, // sfix19_En18 
    input [18:0] Wgt_5_103, // sfix19_En18 
    input [18:0] Wgt_5_104, // sfix19_En18 
    input [18:0] Wgt_5_105, // sfix19_En18 
    input [18:0] Wgt_5_106, // sfix19_En18 
    input [18:0] Wgt_5_107, // sfix19_En18 
    input [18:0] Wgt_5_108, // sfix19_En18 
    input [18:0] Wgt_5_109, // sfix19_En18 
    input [18:0] Wgt_5_110, // sfix19_En18 
    input [18:0] Wgt_5_111, // sfix19_En18 
    input [18:0] Wgt_5_112, // sfix19_En18 
    input [18:0] Wgt_5_113, // sfix19_En18 
    input [18:0] Wgt_5_114, // sfix19_En18 
    input [18:0] Wgt_5_115, // sfix19_En18 
    input [18:0] Wgt_5_116, // sfix19_En18 
    input [18:0] Wgt_5_117, // sfix19_En18 
    input [18:0] Wgt_5_118, // sfix19_En18 
    input [18:0] Wgt_5_119, // sfix19_En18 
    input [18:0] Wgt_5_120, // sfix19_En18 
    input [18:0] Wgt_5_121, // sfix19_En18 
    input [18:0] Wgt_5_122, // sfix19_En18 
    input [18:0] Wgt_5_123, // sfix19_En18 
    input [18:0] Wgt_5_124, // sfix19_En18 
    input [18:0] Wgt_5_125, // sfix19_En18 
    input [18:0] Wgt_5_126, // sfix19_En18 
    input [18:0] Wgt_5_127, // sfix19_En18 
    input [18:0] Wgt_5_128, // sfix19_En18 
    input [18:0] Wgt_5_129, // sfix19_En18 
    input [18:0] Wgt_5_130, // sfix19_En18 
    input [18:0] Wgt_5_131, // sfix19_En18 
    input [18:0] Wgt_5_132, // sfix19_En18 
    input [18:0] Wgt_5_133, // sfix19_En18 
    input [18:0] Wgt_5_134, // sfix19_En18 
    input [18:0] Wgt_5_135, // sfix19_En18 
    input [18:0] Wgt_5_136, // sfix19_En18 
    input [18:0] Wgt_5_137, // sfix19_En18 
    input [18:0] Wgt_5_138, // sfix19_En18 
    input [18:0] Wgt_5_139, // sfix19_En18 
    input [18:0] Wgt_5_140, // sfix19_En18 
    input [18:0] Wgt_5_141, // sfix19_En18 
    input [18:0] Wgt_5_142, // sfix19_En18 
    input [18:0] Wgt_5_143, // sfix19_En18 
    input [18:0] Wgt_5_144, // sfix19_En18 
    input [18:0] Wgt_5_145, // sfix19_En18 
    input [18:0] Wgt_5_146, // sfix19_En18 
    input [18:0] Wgt_5_147, // sfix19_En18 
    input [18:0] Wgt_5_148, // sfix19_En18 
    input [18:0] Wgt_5_149, // sfix19_En18 
    input [18:0] Wgt_5_150, // sfix19_En18 
    input [18:0] Wgt_5_151, // sfix19_En18 
    input [18:0] Wgt_5_152, // sfix19_En18 
    input [18:0] Wgt_5_153, // sfix19_En18 
    input [18:0] Wgt_5_154, // sfix19_En18 
    input [18:0] Wgt_5_155, // sfix19_En18 
    input [18:0] Wgt_5_156, // sfix19_En18 
    input [18:0] Wgt_5_157, // sfix19_En18 
    input [18:0] Wgt_5_158, // sfix19_En18 
    input [18:0] Wgt_5_159, // sfix19_En18 
    input [18:0] Wgt_5_160, // sfix19_En18 
    input [18:0] Wgt_5_161, // sfix19_En18 
    input [18:0] Wgt_5_162, // sfix19_En18 
    input [18:0] Wgt_5_163, // sfix19_En18 
    input [18:0] Wgt_5_164, // sfix19_En18 
    input [18:0] Wgt_5_165, // sfix19_En18 
    input [18:0] Wgt_5_166, // sfix19_En18 
    input [18:0] Wgt_5_167, // sfix19_En18 
    input [18:0] Wgt_5_168, // sfix19_En18 
    input [18:0] Wgt_5_169, // sfix19_En18 
    input [18:0] Wgt_5_170, // sfix19_En18 
    input [18:0] Wgt_5_171, // sfix19_En18 
    input [18:0] Wgt_5_172, // sfix19_En18 
    input [18:0] Wgt_5_173, // sfix19_En18 
    input [18:0] Wgt_5_174, // sfix19_En18 
    input [18:0] Wgt_5_175, // sfix19_En18 
    input [18:0] Wgt_5_176, // sfix19_En18 
    input [18:0] Wgt_5_177, // sfix19_En18 
    input [18:0] Wgt_5_178, // sfix19_En18 
    input [18:0] Wgt_5_179, // sfix19_En18 
    input [18:0] Wgt_5_180, // sfix19_En18 
    input [18:0] Wgt_5_181, // sfix19_En18 
    input [18:0] Wgt_5_182, // sfix19_En18 
    input [18:0] Wgt_5_183, // sfix19_En18 
    input [18:0] Wgt_5_184, // sfix19_En18 
    input [18:0] Wgt_5_185, // sfix19_En18 
    input [18:0] Wgt_5_186, // sfix19_En18 
    input [18:0] Wgt_5_187, // sfix19_En18 
    input [18:0] Wgt_5_188, // sfix19_En18 
    input [18:0] Wgt_5_189, // sfix19_En18 
    input [18:0] Wgt_5_190, // sfix19_En18 
    input [18:0] Wgt_5_191, // sfix19_En18 
    input [18:0] Wgt_5_192, // sfix19_En18 
    input [18:0] Wgt_5_193, // sfix19_En18 
    input [18:0] Wgt_5_194, // sfix19_En18 
    input [18:0] Wgt_5_195, // sfix19_En18 
    input [18:0] Wgt_5_196, // sfix19_En18 
    input [18:0] Wgt_5_197, // sfix19_En18 
    input [18:0] Wgt_5_198, // sfix19_En18 
    input [18:0] Wgt_5_199, // sfix19_En18 
    input [18:0] Wgt_5_200, // sfix19_En18 
    input [18:0] Wgt_5_201, // sfix19_En18 
    input [18:0] Wgt_5_202, // sfix19_En18 
    input [18:0] Wgt_5_203, // sfix19_En18 
    input [18:0] Wgt_5_204, // sfix19_En18 
    input [18:0] Wgt_5_205, // sfix19_En18 
    input [18:0] Wgt_5_206, // sfix19_En18 
    input [18:0] Wgt_5_207, // sfix19_En18 
    input [18:0] Wgt_5_208, // sfix19_En18 
    input [18:0] Wgt_5_209, // sfix19_En18 
    input [18:0] Wgt_5_210, // sfix19_En18 
    input [18:0] Wgt_5_211, // sfix19_En18 
    input [18:0] Wgt_5_212, // sfix19_En18 
    input [18:0] Wgt_5_213, // sfix19_En18 
    input [18:0] Wgt_5_214, // sfix19_En18 
    input [18:0] Wgt_5_215, // sfix19_En18 
    input [18:0] Wgt_5_216, // sfix19_En18 
    input [18:0] Wgt_5_217, // sfix19_En18 
    input [18:0] Wgt_5_218, // sfix19_En18 
    input [18:0] Wgt_5_219, // sfix19_En18 
    input [18:0] Wgt_5_220, // sfix19_En18 
    input [18:0] Wgt_5_221, // sfix19_En18 
    input [18:0] Wgt_5_222, // sfix19_En18 
    input [18:0] Wgt_5_223, // sfix19_En18 
    input [18:0] Wgt_5_224, // sfix19_En18 
    input [18:0] Wgt_5_225, // sfix19_En18 
    input [18:0] Wgt_5_226, // sfix19_En18 
    input [18:0] Wgt_5_227, // sfix19_En18 
    input [18:0] Wgt_5_228, // sfix19_En18 
    input [18:0] Wgt_5_229, // sfix19_En18 
    input [18:0] Wgt_5_230, // sfix19_En18 
    input [18:0] Wgt_5_231, // sfix19_En18 
    input [18:0] Wgt_5_232, // sfix19_En18 
    input [18:0] Wgt_5_233, // sfix19_En18 
    input [18:0] Wgt_5_234, // sfix19_En18 
    input [18:0] Wgt_5_235, // sfix19_En18 
    input [18:0] Wgt_5_236, // sfix19_En18 
    input [18:0] Wgt_5_237, // sfix19_En18 
    input [18:0] Wgt_5_238, // sfix19_En18 
    input [18:0] Wgt_5_239, // sfix19_En18 
    input [18:0] Wgt_5_240, // sfix19_En18 
    input [18:0] Wgt_5_241, // sfix19_En18 
    input [18:0] Wgt_5_242, // sfix19_En18 
    input [18:0] Wgt_5_243, // sfix19_En18 
    input [18:0] Wgt_5_244, // sfix19_En18 
    input [18:0] Wgt_5_245, // sfix19_En18 
    input [18:0] Wgt_5_246, // sfix19_En18 
    input [18:0] Wgt_5_247, // sfix19_En18 
    input [18:0] Wgt_5_248, // sfix19_En18 
    input [18:0] Wgt_5_249, // sfix19_En18 
    input [18:0] Wgt_5_250, // sfix19_En18 
    input [18:0] Wgt_5_251, // sfix19_En18 
    input [18:0] Wgt_5_252, // sfix19_En18 
    input [18:0] Wgt_5_253, // sfix19_En18 
    input [18:0] Wgt_5_254, // sfix19_En18 
    input [18:0] Wgt_5_255, // sfix19_En18 
    input [18:0] Wgt_5_256, // sfix19_En18 
    input [18:0] Wgt_5_257, // sfix19_En18 
    input [18:0] Wgt_5_258, // sfix19_En18 
    input [18:0] Wgt_5_259, // sfix19_En18 
    input [18:0] Wgt_5_260, // sfix19_En18 
    input [18:0] Wgt_5_261, // sfix19_En18 
    input [18:0] Wgt_5_262, // sfix19_En18 
    input [18:0] Wgt_5_263, // sfix19_En18 
    input [18:0] Wgt_5_264, // sfix19_En18 
    input [18:0] Wgt_5_265, // sfix19_En18 
    input [18:0] Wgt_5_266, // sfix19_En18 
    input [18:0] Wgt_5_267, // sfix19_En18 
    input [18:0] Wgt_5_268, // sfix19_En18 
    input [18:0] Wgt_5_269, // sfix19_En18 
    input [18:0] Wgt_5_270, // sfix19_En18 
    input [18:0] Wgt_5_271, // sfix19_En18 
    input [18:0] Wgt_5_272, // sfix19_En18 
    input [18:0] Wgt_5_273, // sfix19_En18 
    input [18:0] Wgt_5_274, // sfix19_En18 
    input [18:0] Wgt_5_275, // sfix19_En18 
    input [18:0] Wgt_5_276, // sfix19_En18 
    input [18:0] Wgt_5_277, // sfix19_En18 
    input [18:0] Wgt_5_278, // sfix19_En18 
    input [18:0] Wgt_5_279, // sfix19_En18 
    input [18:0] Wgt_5_280, // sfix19_En18 
    input [18:0] Wgt_5_281, // sfix19_En18 
    input [18:0] Wgt_5_282, // sfix19_En18 
    input [18:0] Wgt_5_283, // sfix19_En18 
    input [18:0] Wgt_5_284, // sfix19_En18 
    input [18:0] Wgt_5_285, // sfix19_En18 
    input [18:0] Wgt_5_286, // sfix19_En18 
    input [18:0] Wgt_5_287, // sfix19_En18 
    input [18:0] Wgt_5_288, // sfix19_En18 
    input [18:0] Wgt_5_289, // sfix19_En18 
    input [18:0] Wgt_5_290, // sfix19_En18 
    input [18:0] Wgt_5_291, // sfix19_En18 
    input [18:0] Wgt_5_292, // sfix19_En18 
    input [18:0] Wgt_5_293, // sfix19_En18 
    input [18:0] Wgt_5_294, // sfix19_En18 
    input [18:0] Wgt_5_295, // sfix19_En18 
    input [18:0] Wgt_5_296, // sfix19_En18 
    input [18:0] Wgt_5_297, // sfix19_En18 
    input [18:0] Wgt_5_298, // sfix19_En18 
    input [18:0] Wgt_5_299, // sfix19_En18 
    input [18:0] Wgt_5_300, // sfix19_En18 
    input [18:0] Wgt_5_301, // sfix19_En18 
    input [18:0] Wgt_5_302, // sfix19_En18 
    input [18:0] Wgt_5_303, // sfix19_En18 
    input [18:0] Wgt_5_304, // sfix19_En18 
    input [18:0] Wgt_5_305, // sfix19_En18 
    input [18:0] Wgt_5_306, // sfix19_En18 
    input [18:0] Wgt_5_307, // sfix19_En18 
    input [18:0] Wgt_5_308, // sfix19_En18 
    input [18:0] Wgt_5_309, // sfix19_En18 
    input [18:0] Wgt_5_310, // sfix19_En18 
    input [18:0] Wgt_5_311, // sfix19_En18 
    input [18:0] Wgt_5_312, // sfix19_En18 
    input [18:0] Wgt_5_313, // sfix19_En18 
    input [18:0] Wgt_5_314, // sfix19_En18 
    input [18:0] Wgt_5_315, // sfix19_En18 
    input [18:0] Wgt_5_316, // sfix19_En18 
    input [18:0] Wgt_5_317, // sfix19_En18 
    input [18:0] Wgt_5_318, // sfix19_En18 
    input [18:0] Wgt_5_319, // sfix19_En18 
    input [18:0] Wgt_5_320, // sfix19_En18 
    input [18:0] Wgt_5_321, // sfix19_En18 
    input [18:0] Wgt_5_322, // sfix19_En18 
    input [18:0] Wgt_5_323, // sfix19_En18 
    input [18:0] Wgt_5_324, // sfix19_En18 
    input [18:0] Wgt_5_325, // sfix19_En18 
    input [18:0] Wgt_5_326, // sfix19_En18 
    input [18:0] Wgt_5_327, // sfix19_En18 
    input [18:0] Wgt_5_328, // sfix19_En18 
    input [18:0] Wgt_5_329, // sfix19_En18 
    input [18:0] Wgt_5_330, // sfix19_En18 
    input [18:0] Wgt_5_331, // sfix19_En18 
    input [18:0] Wgt_5_332, // sfix19_En18 
    input [18:0] Wgt_5_333, // sfix19_En18 
    input [18:0] Wgt_5_334, // sfix19_En18 
    input [18:0] Wgt_5_335, // sfix19_En18 
    input [18:0] Wgt_5_336, // sfix19_En18 
    input [18:0] Wgt_5_337, // sfix19_En18 
    input [18:0] Wgt_5_338, // sfix19_En18 
    input [18:0] Wgt_5_339, // sfix19_En18 
    input [18:0] Wgt_5_340, // sfix19_En18 
    input [18:0] Wgt_5_341, // sfix19_En18 
    input [18:0] Wgt_5_342, // sfix19_En18 
    input [18:0] Wgt_5_343, // sfix19_En18 
    input [18:0] Wgt_5_344, // sfix19_En18 
    input [18:0] Wgt_5_345, // sfix19_En18 
    input [18:0] Wgt_5_346, // sfix19_En18 
    input [18:0] Wgt_5_347, // sfix19_En18 
    input [18:0] Wgt_5_348, // sfix19_En18 
    input [18:0] Wgt_5_349, // sfix19_En18 
    input [18:0] Wgt_5_350, // sfix19_En18 
    input [18:0] Wgt_5_351, // sfix19_En18 
    input [18:0] Wgt_5_352, // sfix19_En18 
    input [18:0] Wgt_5_353, // sfix19_En18 
    input [18:0] Wgt_5_354, // sfix19_En18 
    input [18:0] Wgt_5_355, // sfix19_En18 
    input [18:0] Wgt_5_356, // sfix19_En18 
    input [18:0] Wgt_5_357, // sfix19_En18 
    input [18:0] Wgt_5_358, // sfix19_En18 
    input [18:0] Wgt_5_359, // sfix19_En18 
    input [18:0] Wgt_5_360, // sfix19_En18 
    input [18:0] Wgt_5_361, // sfix19_En18 
    input [18:0] Wgt_5_362, // sfix19_En18 
    input [18:0] Wgt_5_363, // sfix19_En18 
    input [18:0] Wgt_5_364, // sfix19_En18 
    input [18:0] Wgt_5_365, // sfix19_En18 
    input [18:0] Wgt_5_366, // sfix19_En18 
    input [18:0] Wgt_5_367, // sfix19_En18 
    input [18:0] Wgt_5_368, // sfix19_En18 
    input [18:0] Wgt_5_369, // sfix19_En18 
    input [18:0] Wgt_5_370, // sfix19_En18 
    input [18:0] Wgt_5_371, // sfix19_En18 
    input [18:0] Wgt_5_372, // sfix19_En18 
    input [18:0] Wgt_5_373, // sfix19_En18 
    input [18:0] Wgt_5_374, // sfix19_En18 
    input [18:0] Wgt_5_375, // sfix19_En18 
    input [18:0] Wgt_5_376, // sfix19_En18 
    input [18:0] Wgt_5_377, // sfix19_En18 
    input [18:0] Wgt_5_378, // sfix19_En18 
    input [18:0] Wgt_5_379, // sfix19_En18 
    input [18:0] Wgt_5_380, // sfix19_En18 
    input [18:0] Wgt_5_381, // sfix19_En18 
    input [18:0] Wgt_5_382, // sfix19_En18 
    input [18:0] Wgt_5_383, // sfix19_En18 
    input [18:0] Wgt_5_384, // sfix19_En18 
    input [18:0] Wgt_5_385, // sfix19_En18 
    input [18:0] Wgt_5_386, // sfix19_En18 
    input [18:0] Wgt_5_387, // sfix19_En18 
    input [18:0] Wgt_5_388, // sfix19_En18 
    input [18:0] Wgt_5_389, // sfix19_En18 
    input [18:0] Wgt_5_390, // sfix19_En18 
    input [18:0] Wgt_5_391, // sfix19_En18 
    input [18:0] Wgt_5_392, // sfix19_En18 
    input [18:0] Wgt_5_393, // sfix19_En18 
    input [18:0] Wgt_5_394, // sfix19_En18 
    input [18:0] Wgt_5_395, // sfix19_En18 
    input [18:0] Wgt_5_396, // sfix19_En18 
    input [18:0] Wgt_5_397, // sfix19_En18 
    input [18:0] Wgt_5_398, // sfix19_En18 
    input [18:0] Wgt_5_399, // sfix19_En18 
    input [18:0] Wgt_5_400, // sfix19_En18 
    input [18:0] Wgt_5_401, // sfix19_En18 
    input [18:0] Wgt_5_402, // sfix19_En18 
    input [18:0] Wgt_5_403, // sfix19_En18 
    input [18:0] Wgt_5_404, // sfix19_En18 
    input [18:0] Wgt_5_405, // sfix19_En18 
    input [18:0] Wgt_5_406, // sfix19_En18 
    input [18:0] Wgt_5_407, // sfix19_En18 
    input [18:0] Wgt_5_408, // sfix19_En18 
    input [18:0] Wgt_5_409, // sfix19_En18 
    input [18:0] Wgt_5_410, // sfix19_En18 
    input [18:0] Wgt_5_411, // sfix19_En18 
    input [18:0] Wgt_5_412, // sfix19_En18 
    input [18:0] Wgt_5_413, // sfix19_En18 
    input [18:0] Wgt_5_414, // sfix19_En18 
    input [18:0] Wgt_5_415, // sfix19_En18 
    input [18:0] Wgt_5_416, // sfix19_En18 
    input [18:0] Wgt_5_417, // sfix19_En18 
    input [18:0] Wgt_5_418, // sfix19_En18 
    input [18:0] Wgt_5_419, // sfix19_En18 
    input [18:0] Wgt_5_420, // sfix19_En18 
    input [18:0] Wgt_5_421, // sfix19_En18 
    input [18:0] Wgt_5_422, // sfix19_En18 
    input [18:0] Wgt_5_423, // sfix19_En18 
    input [18:0] Wgt_5_424, // sfix19_En18 
    input [18:0] Wgt_5_425, // sfix19_En18 
    input [18:0] Wgt_5_426, // sfix19_En18 
    input [18:0] Wgt_5_427, // sfix19_En18 
    input [18:0] Wgt_5_428, // sfix19_En18 
    input [18:0] Wgt_5_429, // sfix19_En18 
    input [18:0] Wgt_5_430, // sfix19_En18 
    input [18:0] Wgt_5_431, // sfix19_En18 
    input [18:0] Wgt_5_432, // sfix19_En18 
    input [18:0] Wgt_5_433, // sfix19_En18 
    input [18:0] Wgt_5_434, // sfix19_En18 
    input [18:0] Wgt_5_435, // sfix19_En18 
    input [18:0] Wgt_5_436, // sfix19_En18 
    input [18:0] Wgt_5_437, // sfix19_En18 
    input [18:0] Wgt_5_438, // sfix19_En18 
    input [18:0] Wgt_5_439, // sfix19_En18 
    input [18:0] Wgt_5_440, // sfix19_En18 
    input [18:0] Wgt_5_441, // sfix19_En18 
    input [18:0] Wgt_5_442, // sfix19_En18 
    input [18:0] Wgt_5_443, // sfix19_En18 
    input [18:0] Wgt_5_444, // sfix19_En18 
    input [18:0] Wgt_5_445, // sfix19_En18 
    input [18:0] Wgt_5_446, // sfix19_En18 
    input [18:0] Wgt_5_447, // sfix19_En18 
    input [18:0] Wgt_5_448, // sfix19_En18 
    input [18:0] Wgt_5_449, // sfix19_En18 
    input [18:0] Wgt_5_450, // sfix19_En18 
    input [18:0] Wgt_5_451, // sfix19_En18 
    input [18:0] Wgt_5_452, // sfix19_En18 
    input [18:0] Wgt_5_453, // sfix19_En18 
    input [18:0] Wgt_5_454, // sfix19_En18 
    input [18:0] Wgt_5_455, // sfix19_En18 
    input [18:0] Wgt_5_456, // sfix19_En18 
    input [18:0] Wgt_5_457, // sfix19_En18 
    input [18:0] Wgt_5_458, // sfix19_En18 
    input [18:0] Wgt_5_459, // sfix19_En18 
    input [18:0] Wgt_5_460, // sfix19_En18 
    input [18:0] Wgt_5_461, // sfix19_En18 
    input [18:0] Wgt_5_462, // sfix19_En18 
    input [18:0] Wgt_5_463, // sfix19_En18 
    input [18:0] Wgt_5_464, // sfix19_En18 
    input [18:0] Wgt_5_465, // sfix19_En18 
    input [18:0] Wgt_5_466, // sfix19_En18 
    input [18:0] Wgt_5_467, // sfix19_En18 
    input [18:0] Wgt_5_468, // sfix19_En18 
    input [18:0] Wgt_5_469, // sfix19_En18 
    input [18:0] Wgt_5_470, // sfix19_En18 
    input [18:0] Wgt_5_471, // sfix19_En18 
    input [18:0] Wgt_5_472, // sfix19_En18 
    input [18:0] Wgt_5_473, // sfix19_En18 
    input [18:0] Wgt_5_474, // sfix19_En18 
    input [18:0] Wgt_5_475, // sfix19_En18 
    input [18:0] Wgt_5_476, // sfix19_En18 
    input [18:0] Wgt_5_477, // sfix19_En18 
    input [18:0] Wgt_5_478, // sfix19_En18 
    input [18:0] Wgt_5_479, // sfix19_En18 
    input [18:0] Wgt_5_480, // sfix19_En18 
    input [18:0] Wgt_5_481, // sfix19_En18 
    input [18:0] Wgt_5_482, // sfix19_En18 
    input [18:0] Wgt_5_483, // sfix19_En18 
    input [18:0] Wgt_5_484, // sfix19_En18 
    input [18:0] Wgt_5_485, // sfix19_En18 
    input [18:0] Wgt_5_486, // sfix19_En18 
    input [18:0] Wgt_5_487, // sfix19_En18 
    input [18:0] Wgt_5_488, // sfix19_En18 
    input [18:0] Wgt_5_489, // sfix19_En18 
    input [18:0] Wgt_5_490, // sfix19_En18 
    input [18:0] Wgt_5_491, // sfix19_En18 
    input [18:0] Wgt_5_492, // sfix19_En18 
    input [18:0] Wgt_5_493, // sfix19_En18 
    input [18:0] Wgt_5_494, // sfix19_En18 
    input [18:0] Wgt_5_495, // sfix19_En18 
    input [18:0] Wgt_5_496, // sfix19_En18 
    input [18:0] Wgt_5_497, // sfix19_En18 
    input [18:0] Wgt_5_498, // sfix19_En18 
    input [18:0] Wgt_5_499, // sfix19_En18 
    input [18:0] Wgt_5_500, // sfix19_En18 
    input [18:0] Wgt_5_501, // sfix19_En18 
    input [18:0] Wgt_5_502, // sfix19_En18 
    input [18:0] Wgt_5_503, // sfix19_En18 
    input [18:0] Wgt_5_504, // sfix19_En18 
    input [18:0] Wgt_5_505, // sfix19_En18 
    input [18:0] Wgt_5_506, // sfix19_En18 
    input [18:0] Wgt_5_507, // sfix19_En18 
    input [18:0] Wgt_5_508, // sfix19_En18 
    input [18:0] Wgt_5_509, // sfix19_En18 
    input [18:0] Wgt_5_510, // sfix19_En18 
    input [18:0] Wgt_5_511, // sfix19_En18 
    input [18:0] Wgt_5_512, // sfix19_En18 
    input [18:0] Wgt_5_513, // sfix19_En18 
    input [18:0] Wgt_5_514, // sfix19_En18 
    input [18:0] Wgt_5_515, // sfix19_En18 
    input [18:0] Wgt_5_516, // sfix19_En18 
    input [18:0] Wgt_5_517, // sfix19_En18 
    input [18:0] Wgt_5_518, // sfix19_En18 
    input [18:0] Wgt_5_519, // sfix19_En18 
    input [18:0] Wgt_5_520, // sfix19_En18 
    input [18:0] Wgt_5_521, // sfix19_En18 
    input [18:0] Wgt_5_522, // sfix19_En18 
    input [18:0] Wgt_5_523, // sfix19_En18 
    input [18:0] Wgt_5_524, // sfix19_En18 
    input [18:0] Wgt_5_525, // sfix19_En18 
    input [18:0] Wgt_5_526, // sfix19_En18 
    input [18:0] Wgt_5_527, // sfix19_En18 
    input [18:0] Wgt_5_528, // sfix19_En18 
    input [18:0] Wgt_5_529, // sfix19_En18 
    input [18:0] Wgt_5_530, // sfix19_En18 
    input [18:0] Wgt_5_531, // sfix19_En18 
    input [18:0] Wgt_5_532, // sfix19_En18 
    input [18:0] Wgt_5_533, // sfix19_En18 
    input [18:0] Wgt_5_534, // sfix19_En18 
    input [18:0] Wgt_5_535, // sfix19_En18 
    input [18:0] Wgt_5_536, // sfix19_En18 
    input [18:0] Wgt_5_537, // sfix19_En18 
    input [18:0] Wgt_5_538, // sfix19_En18 
    input [18:0] Wgt_5_539, // sfix19_En18 
    input [18:0] Wgt_5_540, // sfix19_En18 
    input [18:0] Wgt_5_541, // sfix19_En18 
    input [18:0] Wgt_5_542, // sfix19_En18 
    input [18:0] Wgt_5_543, // sfix19_En18 
    input [18:0] Wgt_5_544, // sfix19_En18 
    input [18:0] Wgt_5_545, // sfix19_En18 
    input [18:0] Wgt_5_546, // sfix19_En18 
    input [18:0] Wgt_5_547, // sfix19_En18 
    input [18:0] Wgt_5_548, // sfix19_En18 
    input [18:0] Wgt_5_549, // sfix19_En18 
    input [18:0] Wgt_5_550, // sfix19_En18 
    input [18:0] Wgt_5_551, // sfix19_En18 
    input [18:0] Wgt_5_552, // sfix19_En18 
    input [18:0] Wgt_5_553, // sfix19_En18 
    input [18:0] Wgt_5_554, // sfix19_En18 
    input [18:0] Wgt_5_555, // sfix19_En18 
    input [18:0] Wgt_5_556, // sfix19_En18 
    input [18:0] Wgt_5_557, // sfix19_En18 
    input [18:0] Wgt_5_558, // sfix19_En18 
    input [18:0] Wgt_5_559, // sfix19_En18 
    input [18:0] Wgt_5_560, // sfix19_En18 
    input [18:0] Wgt_5_561, // sfix19_En18 
    input [18:0] Wgt_5_562, // sfix19_En18 
    input [18:0] Wgt_5_563, // sfix19_En18 
    input [18:0] Wgt_5_564, // sfix19_En18 
    input [18:0] Wgt_5_565, // sfix19_En18 
    input [18:0] Wgt_5_566, // sfix19_En18 
    input [18:0] Wgt_5_567, // sfix19_En18 
    input [18:0] Wgt_5_568, // sfix19_En18 
    input [18:0] Wgt_5_569, // sfix19_En18 
    input [18:0] Wgt_5_570, // sfix19_En18 
    input [18:0] Wgt_5_571, // sfix19_En18 
    input [18:0] Wgt_5_572, // sfix19_En18 
    input [18:0] Wgt_5_573, // sfix19_En18 
    input [18:0] Wgt_5_574, // sfix19_En18 
    input [18:0] Wgt_5_575, // sfix19_En18 
    input [18:0] Wgt_5_576, // sfix19_En18 
    input [18:0] Wgt_5_577, // sfix19_En18 
    input [18:0] Wgt_5_578, // sfix19_En18 
    input [18:0] Wgt_5_579, // sfix19_En18 
    input [18:0] Wgt_5_580, // sfix19_En18 
    input [18:0] Wgt_5_581, // sfix19_En18 
    input [18:0] Wgt_5_582, // sfix19_En18 
    input [18:0] Wgt_5_583, // sfix19_En18 
    input [18:0] Wgt_5_584, // sfix19_En18 
    input [18:0] Wgt_5_585, // sfix19_En18 
    input [18:0] Wgt_5_586, // sfix19_En18 
    input [18:0] Wgt_5_587, // sfix19_En18 
    input [18:0] Wgt_5_588, // sfix19_En18 
    input [18:0] Wgt_5_589, // sfix19_En18 
    input [18:0] Wgt_5_590, // sfix19_En18 
    input [18:0] Wgt_5_591, // sfix19_En18 
    input [18:0] Wgt_5_592, // sfix19_En18 
    input [18:0] Wgt_5_593, // sfix19_En18 
    input [18:0] Wgt_5_594, // sfix19_En18 
    input [18:0] Wgt_5_595, // sfix19_En18 
    input [18:0] Wgt_5_596, // sfix19_En18 
    input [18:0] Wgt_5_597, // sfix19_En18 
    input [18:0] Wgt_5_598, // sfix19_En18 
    input [18:0] Wgt_5_599, // sfix19_En18 
    input [18:0] Wgt_5_600, // sfix19_En18 
    input [18:0] Wgt_5_601, // sfix19_En18 
    input [18:0] Wgt_5_602, // sfix19_En18 
    input [18:0] Wgt_5_603, // sfix19_En18 
    input [18:0] Wgt_5_604, // sfix19_En18 
    input [18:0] Wgt_5_605, // sfix19_En18 
    input [18:0] Wgt_5_606, // sfix19_En18 
    input [18:0] Wgt_5_607, // sfix19_En18 
    input [18:0] Wgt_5_608, // sfix19_En18 
    input [18:0] Wgt_5_609, // sfix19_En18 
    input [18:0] Wgt_5_610, // sfix19_En18 
    input [18:0] Wgt_5_611, // sfix19_En18 
    input [18:0] Wgt_5_612, // sfix19_En18 
    input [18:0] Wgt_5_613, // sfix19_En18 
    input [18:0] Wgt_5_614, // sfix19_En18 
    input [18:0] Wgt_5_615, // sfix19_En18 
    input [18:0] Wgt_5_616, // sfix19_En18 
    input [18:0] Wgt_5_617, // sfix19_En18 
    input [18:0] Wgt_5_618, // sfix19_En18 
    input [18:0] Wgt_5_619, // sfix19_En18 
    input [18:0] Wgt_5_620, // sfix19_En18 
    input [18:0] Wgt_5_621, // sfix19_En18 
    input [18:0] Wgt_5_622, // sfix19_En18 
    input [18:0] Wgt_5_623, // sfix19_En18 
    input [18:0] Wgt_5_624, // sfix19_En18 
    input [18:0] Wgt_5_625, // sfix19_En18 
    input [18:0] Wgt_5_626, // sfix19_En18 
    input [18:0] Wgt_5_627, // sfix19_En18 
    input [18:0] Wgt_5_628, // sfix19_En18 
    input [18:0] Wgt_5_629, // sfix19_En18 
    input [18:0] Wgt_5_630, // sfix19_En18 
    input [18:0] Wgt_5_631, // sfix19_En18 
    input [18:0] Wgt_5_632, // sfix19_En18 
    input [18:0] Wgt_5_633, // sfix19_En18 
    input [18:0] Wgt_5_634, // sfix19_En18 
    input [18:0] Wgt_5_635, // sfix19_En18 
    input [18:0] Wgt_5_636, // sfix19_En18 
    input [18:0] Wgt_5_637, // sfix19_En18 
    input [18:0] Wgt_5_638, // sfix19_En18 
    input [18:0] Wgt_5_639, // sfix19_En18 
    input [18:0] Wgt_5_640, // sfix19_En18 
    input [18:0] Wgt_5_641, // sfix19_En18 
    input [18:0] Wgt_5_642, // sfix19_En18 
    input [18:0] Wgt_5_643, // sfix19_En18 
    input [18:0] Wgt_5_644, // sfix19_En18 
    input [18:0] Wgt_5_645, // sfix19_En18 
    input [18:0] Wgt_5_646, // sfix19_En18 
    input [18:0] Wgt_5_647, // sfix19_En18 
    input [18:0] Wgt_5_648, // sfix19_En18 
    input [18:0] Wgt_5_649, // sfix19_En18 
    input [18:0] Wgt_5_650, // sfix19_En18 
    input [18:0] Wgt_5_651, // sfix19_En18 
    input [18:0] Wgt_5_652, // sfix19_En18 
    input [18:0] Wgt_5_653, // sfix19_En18 
    input [18:0] Wgt_5_654, // sfix19_En18 
    input [18:0] Wgt_5_655, // sfix19_En18 
    input [18:0] Wgt_5_656, // sfix19_En18 
    input [18:0] Wgt_5_657, // sfix19_En18 
    input [18:0] Wgt_5_658, // sfix19_En18 
    input [18:0] Wgt_5_659, // sfix19_En18 
    input [18:0] Wgt_5_660, // sfix19_En18 
    input [18:0] Wgt_5_661, // sfix19_En18 
    input [18:0] Wgt_5_662, // sfix19_En18 
    input [18:0] Wgt_5_663, // sfix19_En18 
    input [18:0] Wgt_5_664, // sfix19_En18 
    input [18:0] Wgt_5_665, // sfix19_En18 
    input [18:0] Wgt_5_666, // sfix19_En18 
    input [18:0] Wgt_5_667, // sfix19_En18 
    input [18:0] Wgt_5_668, // sfix19_En18 
    input [18:0] Wgt_5_669, // sfix19_En18 
    input [18:0] Wgt_5_670, // sfix19_En18 
    input [18:0] Wgt_5_671, // sfix19_En18 
    input [18:0] Wgt_5_672, // sfix19_En18 
    input [18:0] Wgt_5_673, // sfix19_En18 
    input [18:0] Wgt_5_674, // sfix19_En18 
    input [18:0] Wgt_5_675, // sfix19_En18 
    input [18:0] Wgt_5_676, // sfix19_En18 
    input [18:0] Wgt_5_677, // sfix19_En18 
    input [18:0] Wgt_5_678, // sfix19_En18 
    input [18:0] Wgt_5_679, // sfix19_En18 
    input [18:0] Wgt_5_680, // sfix19_En18 
    input [18:0] Wgt_5_681, // sfix19_En18 
    input [18:0] Wgt_5_682, // sfix19_En18 
    input [18:0] Wgt_5_683, // sfix19_En18 
    input [18:0] Wgt_5_684, // sfix19_En18 
    input [18:0] Wgt_5_685, // sfix19_En18 
    input [18:0] Wgt_5_686, // sfix19_En18 
    input [18:0] Wgt_5_687, // sfix19_En18 
    input [18:0] Wgt_5_688, // sfix19_En18 
    input [18:0] Wgt_5_689, // sfix19_En18 
    input [18:0] Wgt_5_690, // sfix19_En18 
    input [18:0] Wgt_5_691, // sfix19_En18 
    input [18:0] Wgt_5_692, // sfix19_En18 
    input [18:0] Wgt_5_693, // sfix19_En18 
    input [18:0] Wgt_5_694, // sfix19_En18 
    input [18:0] Wgt_5_695, // sfix19_En18 
    input [18:0] Wgt_5_696, // sfix19_En18 
    input [18:0] Wgt_5_697, // sfix19_En18 
    input [18:0] Wgt_5_698, // sfix19_En18 
    input [18:0] Wgt_5_699, // sfix19_En18 
    input [18:0] Wgt_5_700, // sfix19_En18 
    input [18:0] Wgt_5_701, // sfix19_En18 
    input [18:0] Wgt_5_702, // sfix19_En18 
    input [18:0] Wgt_5_703, // sfix19_En18 
    input [18:0] Wgt_5_704, // sfix19_En18 
    input [18:0] Wgt_5_705, // sfix19_En18 
    input [18:0] Wgt_5_706, // sfix19_En18 
    input [18:0] Wgt_5_707, // sfix19_En18 
    input [18:0] Wgt_5_708, // sfix19_En18 
    input [18:0] Wgt_5_709, // sfix19_En18 
    input [18:0] Wgt_5_710, // sfix19_En18 
    input [18:0] Wgt_5_711, // sfix19_En18 
    input [18:0] Wgt_5_712, // sfix19_En18 
    input [18:0] Wgt_5_713, // sfix19_En18 
    input [18:0] Wgt_5_714, // sfix19_En18 
    input [18:0] Wgt_5_715, // sfix19_En18 
    input [18:0] Wgt_5_716, // sfix19_En18 
    input [18:0] Wgt_5_717, // sfix19_En18 
    input [18:0] Wgt_5_718, // sfix19_En18 
    input [18:0] Wgt_5_719, // sfix19_En18 
    input [18:0] Wgt_5_720, // sfix19_En18 
    input [18:0] Wgt_5_721, // sfix19_En18 
    input [18:0] Wgt_5_722, // sfix19_En18 
    input [18:0] Wgt_5_723, // sfix19_En18 
    input [18:0] Wgt_5_724, // sfix19_En18 
    input [18:0] Wgt_5_725, // sfix19_En18 
    input [18:0] Wgt_5_726, // sfix19_En18 
    input [18:0] Wgt_5_727, // sfix19_En18 
    input [18:0] Wgt_5_728, // sfix19_En18 
    input [18:0] Wgt_5_729, // sfix19_En18 
    input [18:0] Wgt_5_730, // sfix19_En18 
    input [18:0] Wgt_5_731, // sfix19_En18 
    input [18:0] Wgt_5_732, // sfix19_En18 
    input [18:0] Wgt_5_733, // sfix19_En18 
    input [18:0] Wgt_5_734, // sfix19_En18 
    input [18:0] Wgt_5_735, // sfix19_En18 
    input [18:0] Wgt_5_736, // sfix19_En18 
    input [18:0] Wgt_5_737, // sfix19_En18 
    input [18:0] Wgt_5_738, // sfix19_En18 
    input [18:0] Wgt_5_739, // sfix19_En18 
    input [18:0] Wgt_5_740, // sfix19_En18 
    input [18:0] Wgt_5_741, // sfix19_En18 
    input [18:0] Wgt_5_742, // sfix19_En18 
    input [18:0] Wgt_5_743, // sfix19_En18 
    input [18:0] Wgt_5_744, // sfix19_En18 
    input [18:0] Wgt_5_745, // sfix19_En18 
    input [18:0] Wgt_5_746, // sfix19_En18 
    input [18:0] Wgt_5_747, // sfix19_En18 
    input [18:0] Wgt_5_748, // sfix19_En18 
    input [18:0] Wgt_5_749, // sfix19_En18 
    input [18:0] Wgt_5_750, // sfix19_En18 
    input [18:0] Wgt_5_751, // sfix19_En18 
    input [18:0] Wgt_5_752, // sfix19_En18 
    input [18:0] Wgt_5_753, // sfix19_En18 
    input [18:0] Wgt_5_754, // sfix19_En18 
    input [18:0] Wgt_5_755, // sfix19_En18 
    input [18:0] Wgt_5_756, // sfix19_En18 
    input [18:0] Wgt_5_757, // sfix19_En18 
    input [18:0] Wgt_5_758, // sfix19_En18 
    input [18:0] Wgt_5_759, // sfix19_En18 
    input [18:0] Wgt_5_760, // sfix19_En18 
    input [18:0] Wgt_5_761, // sfix19_En18 
    input [18:0] Wgt_5_762, // sfix19_En18 
    input [18:0] Wgt_5_763, // sfix19_En18 
    input [18:0] Wgt_5_764, // sfix19_En18 
    input [18:0] Wgt_5_765, // sfix19_En18 
    input [18:0] Wgt_5_766, // sfix19_En18 
    input [18:0] Wgt_5_767, // sfix19_En18 
    input [18:0] Wgt_5_768, // sfix19_En18 
    input [18:0] Wgt_5_769, // sfix19_En18 
    input [18:0] Wgt_5_770, // sfix19_En18 
    input [18:0] Wgt_5_771, // sfix19_En18 
    input [18:0] Wgt_5_772, // sfix19_En18 
    input [18:0] Wgt_5_773, // sfix19_En18 
    input [18:0] Wgt_5_774, // sfix19_En18 
    input [18:0] Wgt_5_775, // sfix19_En18 
    input [18:0] Wgt_5_776, // sfix19_En18 
    input [18:0] Wgt_5_777, // sfix19_En18 
    input [18:0] Wgt_5_778, // sfix19_En18 
    input [18:0] Wgt_5_779, // sfix19_En18 
    input [18:0] Wgt_5_780, // sfix19_En18 
    input [18:0] Wgt_5_781, // sfix19_En18 
    input [18:0] Wgt_5_782, // sfix19_En18 
    input [18:0] Wgt_5_783, // sfix19_En18 
    input [18:0] Wgt_5_784, // sfix19_En18 
    input [18:0] Wgt_6_0, // sfix19_En18 
    input [18:0] Wgt_6_1, // sfix19_En18 
    input [18:0] Wgt_6_2, // sfix19_En18 
    input [18:0] Wgt_6_3, // sfix19_En18 
    input [18:0] Wgt_6_4, // sfix19_En18 
    input [18:0] Wgt_6_5, // sfix19_En18 
    input [18:0] Wgt_6_6, // sfix19_En18 
    input [18:0] Wgt_6_7, // sfix19_En18 
    input [18:0] Wgt_6_8, // sfix19_En18 
    input [18:0] Wgt_6_9, // sfix19_En18 
    input [18:0] Wgt_6_10, // sfix19_En18 
    input [18:0] Wgt_6_11, // sfix19_En18 
    input [18:0] Wgt_6_12, // sfix19_En18 
    input [18:0] Wgt_6_13, // sfix19_En18 
    input [18:0] Wgt_6_14, // sfix19_En18 
    input [18:0] Wgt_6_15, // sfix19_En18 
    input [18:0] Wgt_6_16, // sfix19_En18 
    input [18:0] Wgt_6_17, // sfix19_En18 
    input [18:0] Wgt_6_18, // sfix19_En18 
    input [18:0] Wgt_6_19, // sfix19_En18 
    input [18:0] Wgt_6_20, // sfix19_En18 
    input [18:0] Wgt_6_21, // sfix19_En18 
    input [18:0] Wgt_6_22, // sfix19_En18 
    input [18:0] Wgt_6_23, // sfix19_En18 
    input [18:0] Wgt_6_24, // sfix19_En18 
    input [18:0] Wgt_6_25, // sfix19_En18 
    input [18:0] Wgt_6_26, // sfix19_En18 
    input [18:0] Wgt_6_27, // sfix19_En18 
    input [18:0] Wgt_6_28, // sfix19_En18 
    input [18:0] Wgt_6_29, // sfix19_En18 
    input [18:0] Wgt_6_30, // sfix19_En18 
    input [18:0] Wgt_6_31, // sfix19_En18 
    input [18:0] Wgt_6_32, // sfix19_En18 
    input [18:0] Wgt_6_33, // sfix19_En18 
    input [18:0] Wgt_6_34, // sfix19_En18 
    input [18:0] Wgt_6_35, // sfix19_En18 
    input [18:0] Wgt_6_36, // sfix19_En18 
    input [18:0] Wgt_6_37, // sfix19_En18 
    input [18:0] Wgt_6_38, // sfix19_En18 
    input [18:0] Wgt_6_39, // sfix19_En18 
    input [18:0] Wgt_6_40, // sfix19_En18 
    input [18:0] Wgt_6_41, // sfix19_En18 
    input [18:0] Wgt_6_42, // sfix19_En18 
    input [18:0] Wgt_6_43, // sfix19_En18 
    input [18:0] Wgt_6_44, // sfix19_En18 
    input [18:0] Wgt_6_45, // sfix19_En18 
    input [18:0] Wgt_6_46, // sfix19_En18 
    input [18:0] Wgt_6_47, // sfix19_En18 
    input [18:0] Wgt_6_48, // sfix19_En18 
    input [18:0] Wgt_6_49, // sfix19_En18 
    input [18:0] Wgt_6_50, // sfix19_En18 
    input [18:0] Wgt_6_51, // sfix19_En18 
    input [18:0] Wgt_6_52, // sfix19_En18 
    input [18:0] Wgt_6_53, // sfix19_En18 
    input [18:0] Wgt_6_54, // sfix19_En18 
    input [18:0] Wgt_6_55, // sfix19_En18 
    input [18:0] Wgt_6_56, // sfix19_En18 
    input [18:0] Wgt_6_57, // sfix19_En18 
    input [18:0] Wgt_6_58, // sfix19_En18 
    input [18:0] Wgt_6_59, // sfix19_En18 
    input [18:0] Wgt_6_60, // sfix19_En18 
    input [18:0] Wgt_6_61, // sfix19_En18 
    input [18:0] Wgt_6_62, // sfix19_En18 
    input [18:0] Wgt_6_63, // sfix19_En18 
    input [18:0] Wgt_6_64, // sfix19_En18 
    input [18:0] Wgt_6_65, // sfix19_En18 
    input [18:0] Wgt_6_66, // sfix19_En18 
    input [18:0] Wgt_6_67, // sfix19_En18 
    input [18:0] Wgt_6_68, // sfix19_En18 
    input [18:0] Wgt_6_69, // sfix19_En18 
    input [18:0] Wgt_6_70, // sfix19_En18 
    input [18:0] Wgt_6_71, // sfix19_En18 
    input [18:0] Wgt_6_72, // sfix19_En18 
    input [18:0] Wgt_6_73, // sfix19_En18 
    input [18:0] Wgt_6_74, // sfix19_En18 
    input [18:0] Wgt_6_75, // sfix19_En18 
    input [18:0] Wgt_6_76, // sfix19_En18 
    input [18:0] Wgt_6_77, // sfix19_En18 
    input [18:0] Wgt_6_78, // sfix19_En18 
    input [18:0] Wgt_6_79, // sfix19_En18 
    input [18:0] Wgt_6_80, // sfix19_En18 
    input [18:0] Wgt_6_81, // sfix19_En18 
    input [18:0] Wgt_6_82, // sfix19_En18 
    input [18:0] Wgt_6_83, // sfix19_En18 
    input [18:0] Wgt_6_84, // sfix19_En18 
    input [18:0] Wgt_6_85, // sfix19_En18 
    input [18:0] Wgt_6_86, // sfix19_En18 
    input [18:0] Wgt_6_87, // sfix19_En18 
    input [18:0] Wgt_6_88, // sfix19_En18 
    input [18:0] Wgt_6_89, // sfix19_En18 
    input [18:0] Wgt_6_90, // sfix19_En18 
    input [18:0] Wgt_6_91, // sfix19_En18 
    input [18:0] Wgt_6_92, // sfix19_En18 
    input [18:0] Wgt_6_93, // sfix19_En18 
    input [18:0] Wgt_6_94, // sfix19_En18 
    input [18:0] Wgt_6_95, // sfix19_En18 
    input [18:0] Wgt_6_96, // sfix19_En18 
    input [18:0] Wgt_6_97, // sfix19_En18 
    input [18:0] Wgt_6_98, // sfix19_En18 
    input [18:0] Wgt_6_99, // sfix19_En18 
    input [18:0] Wgt_6_100, // sfix19_En18 
    input [18:0] Wgt_6_101, // sfix19_En18 
    input [18:0] Wgt_6_102, // sfix19_En18 
    input [18:0] Wgt_6_103, // sfix19_En18 
    input [18:0] Wgt_6_104, // sfix19_En18 
    input [18:0] Wgt_6_105, // sfix19_En18 
    input [18:0] Wgt_6_106, // sfix19_En18 
    input [18:0] Wgt_6_107, // sfix19_En18 
    input [18:0] Wgt_6_108, // sfix19_En18 
    input [18:0] Wgt_6_109, // sfix19_En18 
    input [18:0] Wgt_6_110, // sfix19_En18 
    input [18:0] Wgt_6_111, // sfix19_En18 
    input [18:0] Wgt_6_112, // sfix19_En18 
    input [18:0] Wgt_6_113, // sfix19_En18 
    input [18:0] Wgt_6_114, // sfix19_En18 
    input [18:0] Wgt_6_115, // sfix19_En18 
    input [18:0] Wgt_6_116, // sfix19_En18 
    input [18:0] Wgt_6_117, // sfix19_En18 
    input [18:0] Wgt_6_118, // sfix19_En18 
    input [18:0] Wgt_6_119, // sfix19_En18 
    input [18:0] Wgt_6_120, // sfix19_En18 
    input [18:0] Wgt_6_121, // sfix19_En18 
    input [18:0] Wgt_6_122, // sfix19_En18 
    input [18:0] Wgt_6_123, // sfix19_En18 
    input [18:0] Wgt_6_124, // sfix19_En18 
    input [18:0] Wgt_6_125, // sfix19_En18 
    input [18:0] Wgt_6_126, // sfix19_En18 
    input [18:0] Wgt_6_127, // sfix19_En18 
    input [18:0] Wgt_6_128, // sfix19_En18 
    input [18:0] Wgt_6_129, // sfix19_En18 
    input [18:0] Wgt_6_130, // sfix19_En18 
    input [18:0] Wgt_6_131, // sfix19_En18 
    input [18:0] Wgt_6_132, // sfix19_En18 
    input [18:0] Wgt_6_133, // sfix19_En18 
    input [18:0] Wgt_6_134, // sfix19_En18 
    input [18:0] Wgt_6_135, // sfix19_En18 
    input [18:0] Wgt_6_136, // sfix19_En18 
    input [18:0] Wgt_6_137, // sfix19_En18 
    input [18:0] Wgt_6_138, // sfix19_En18 
    input [18:0] Wgt_6_139, // sfix19_En18 
    input [18:0] Wgt_6_140, // sfix19_En18 
    input [18:0] Wgt_6_141, // sfix19_En18 
    input [18:0] Wgt_6_142, // sfix19_En18 
    input [18:0] Wgt_6_143, // sfix19_En18 
    input [18:0] Wgt_6_144, // sfix19_En18 
    input [18:0] Wgt_6_145, // sfix19_En18 
    input [18:0] Wgt_6_146, // sfix19_En18 
    input [18:0] Wgt_6_147, // sfix19_En18 
    input [18:0] Wgt_6_148, // sfix19_En18 
    input [18:0] Wgt_6_149, // sfix19_En18 
    input [18:0] Wgt_6_150, // sfix19_En18 
    input [18:0] Wgt_6_151, // sfix19_En18 
    input [18:0] Wgt_6_152, // sfix19_En18 
    input [18:0] Wgt_6_153, // sfix19_En18 
    input [18:0] Wgt_6_154, // sfix19_En18 
    input [18:0] Wgt_6_155, // sfix19_En18 
    input [18:0] Wgt_6_156, // sfix19_En18 
    input [18:0] Wgt_6_157, // sfix19_En18 
    input [18:0] Wgt_6_158, // sfix19_En18 
    input [18:0] Wgt_6_159, // sfix19_En18 
    input [18:0] Wgt_6_160, // sfix19_En18 
    input [18:0] Wgt_6_161, // sfix19_En18 
    input [18:0] Wgt_6_162, // sfix19_En18 
    input [18:0] Wgt_6_163, // sfix19_En18 
    input [18:0] Wgt_6_164, // sfix19_En18 
    input [18:0] Wgt_6_165, // sfix19_En18 
    input [18:0] Wgt_6_166, // sfix19_En18 
    input [18:0] Wgt_6_167, // sfix19_En18 
    input [18:0] Wgt_6_168, // sfix19_En18 
    input [18:0] Wgt_6_169, // sfix19_En18 
    input [18:0] Wgt_6_170, // sfix19_En18 
    input [18:0] Wgt_6_171, // sfix19_En18 
    input [18:0] Wgt_6_172, // sfix19_En18 
    input [18:0] Wgt_6_173, // sfix19_En18 
    input [18:0] Wgt_6_174, // sfix19_En18 
    input [18:0] Wgt_6_175, // sfix19_En18 
    input [18:0] Wgt_6_176, // sfix19_En18 
    input [18:0] Wgt_6_177, // sfix19_En18 
    input [18:0] Wgt_6_178, // sfix19_En18 
    input [18:0] Wgt_6_179, // sfix19_En18 
    input [18:0] Wgt_6_180, // sfix19_En18 
    input [18:0] Wgt_6_181, // sfix19_En18 
    input [18:0] Wgt_6_182, // sfix19_En18 
    input [18:0] Wgt_6_183, // sfix19_En18 
    input [18:0] Wgt_6_184, // sfix19_En18 
    input [18:0] Wgt_6_185, // sfix19_En18 
    input [18:0] Wgt_6_186, // sfix19_En18 
    input [18:0] Wgt_6_187, // sfix19_En18 
    input [18:0] Wgt_6_188, // sfix19_En18 
    input [18:0] Wgt_6_189, // sfix19_En18 
    input [18:0] Wgt_6_190, // sfix19_En18 
    input [18:0] Wgt_6_191, // sfix19_En18 
    input [18:0] Wgt_6_192, // sfix19_En18 
    input [18:0] Wgt_6_193, // sfix19_En18 
    input [18:0] Wgt_6_194, // sfix19_En18 
    input [18:0] Wgt_6_195, // sfix19_En18 
    input [18:0] Wgt_6_196, // sfix19_En18 
    input [18:0] Wgt_6_197, // sfix19_En18 
    input [18:0] Wgt_6_198, // sfix19_En18 
    input [18:0] Wgt_6_199, // sfix19_En18 
    input [18:0] Wgt_6_200, // sfix19_En18 
    input [18:0] Wgt_6_201, // sfix19_En18 
    input [18:0] Wgt_6_202, // sfix19_En18 
    input [18:0] Wgt_6_203, // sfix19_En18 
    input [18:0] Wgt_6_204, // sfix19_En18 
    input [18:0] Wgt_6_205, // sfix19_En18 
    input [18:0] Wgt_6_206, // sfix19_En18 
    input [18:0] Wgt_6_207, // sfix19_En18 
    input [18:0] Wgt_6_208, // sfix19_En18 
    input [18:0] Wgt_6_209, // sfix19_En18 
    input [18:0] Wgt_6_210, // sfix19_En18 
    input [18:0] Wgt_6_211, // sfix19_En18 
    input [18:0] Wgt_6_212, // sfix19_En18 
    input [18:0] Wgt_6_213, // sfix19_En18 
    input [18:0] Wgt_6_214, // sfix19_En18 
    input [18:0] Wgt_6_215, // sfix19_En18 
    input [18:0] Wgt_6_216, // sfix19_En18 
    input [18:0] Wgt_6_217, // sfix19_En18 
    input [18:0] Wgt_6_218, // sfix19_En18 
    input [18:0] Wgt_6_219, // sfix19_En18 
    input [18:0] Wgt_6_220, // sfix19_En18 
    input [18:0] Wgt_6_221, // sfix19_En18 
    input [18:0] Wgt_6_222, // sfix19_En18 
    input [18:0] Wgt_6_223, // sfix19_En18 
    input [18:0] Wgt_6_224, // sfix19_En18 
    input [18:0] Wgt_6_225, // sfix19_En18 
    input [18:0] Wgt_6_226, // sfix19_En18 
    input [18:0] Wgt_6_227, // sfix19_En18 
    input [18:0] Wgt_6_228, // sfix19_En18 
    input [18:0] Wgt_6_229, // sfix19_En18 
    input [18:0] Wgt_6_230, // sfix19_En18 
    input [18:0] Wgt_6_231, // sfix19_En18 
    input [18:0] Wgt_6_232, // sfix19_En18 
    input [18:0] Wgt_6_233, // sfix19_En18 
    input [18:0] Wgt_6_234, // sfix19_En18 
    input [18:0] Wgt_6_235, // sfix19_En18 
    input [18:0] Wgt_6_236, // sfix19_En18 
    input [18:0] Wgt_6_237, // sfix19_En18 
    input [18:0] Wgt_6_238, // sfix19_En18 
    input [18:0] Wgt_6_239, // sfix19_En18 
    input [18:0] Wgt_6_240, // sfix19_En18 
    input [18:0] Wgt_6_241, // sfix19_En18 
    input [18:0] Wgt_6_242, // sfix19_En18 
    input [18:0] Wgt_6_243, // sfix19_En18 
    input [18:0] Wgt_6_244, // sfix19_En18 
    input [18:0] Wgt_6_245, // sfix19_En18 
    input [18:0] Wgt_6_246, // sfix19_En18 
    input [18:0] Wgt_6_247, // sfix19_En18 
    input [18:0] Wgt_6_248, // sfix19_En18 
    input [18:0] Wgt_6_249, // sfix19_En18 
    input [18:0] Wgt_6_250, // sfix19_En18 
    input [18:0] Wgt_6_251, // sfix19_En18 
    input [18:0] Wgt_6_252, // sfix19_En18 
    input [18:0] Wgt_6_253, // sfix19_En18 
    input [18:0] Wgt_6_254, // sfix19_En18 
    input [18:0] Wgt_6_255, // sfix19_En18 
    input [18:0] Wgt_6_256, // sfix19_En18 
    input [18:0] Wgt_6_257, // sfix19_En18 
    input [18:0] Wgt_6_258, // sfix19_En18 
    input [18:0] Wgt_6_259, // sfix19_En18 
    input [18:0] Wgt_6_260, // sfix19_En18 
    input [18:0] Wgt_6_261, // sfix19_En18 
    input [18:0] Wgt_6_262, // sfix19_En18 
    input [18:0] Wgt_6_263, // sfix19_En18 
    input [18:0] Wgt_6_264, // sfix19_En18 
    input [18:0] Wgt_6_265, // sfix19_En18 
    input [18:0] Wgt_6_266, // sfix19_En18 
    input [18:0] Wgt_6_267, // sfix19_En18 
    input [18:0] Wgt_6_268, // sfix19_En18 
    input [18:0] Wgt_6_269, // sfix19_En18 
    input [18:0] Wgt_6_270, // sfix19_En18 
    input [18:0] Wgt_6_271, // sfix19_En18 
    input [18:0] Wgt_6_272, // sfix19_En18 
    input [18:0] Wgt_6_273, // sfix19_En18 
    input [18:0] Wgt_6_274, // sfix19_En18 
    input [18:0] Wgt_6_275, // sfix19_En18 
    input [18:0] Wgt_6_276, // sfix19_En18 
    input [18:0] Wgt_6_277, // sfix19_En18 
    input [18:0] Wgt_6_278, // sfix19_En18 
    input [18:0] Wgt_6_279, // sfix19_En18 
    input [18:0] Wgt_6_280, // sfix19_En18 
    input [18:0] Wgt_6_281, // sfix19_En18 
    input [18:0] Wgt_6_282, // sfix19_En18 
    input [18:0] Wgt_6_283, // sfix19_En18 
    input [18:0] Wgt_6_284, // sfix19_En18 
    input [18:0] Wgt_6_285, // sfix19_En18 
    input [18:0] Wgt_6_286, // sfix19_En18 
    input [18:0] Wgt_6_287, // sfix19_En18 
    input [18:0] Wgt_6_288, // sfix19_En18 
    input [18:0] Wgt_6_289, // sfix19_En18 
    input [18:0] Wgt_6_290, // sfix19_En18 
    input [18:0] Wgt_6_291, // sfix19_En18 
    input [18:0] Wgt_6_292, // sfix19_En18 
    input [18:0] Wgt_6_293, // sfix19_En18 
    input [18:0] Wgt_6_294, // sfix19_En18 
    input [18:0] Wgt_6_295, // sfix19_En18 
    input [18:0] Wgt_6_296, // sfix19_En18 
    input [18:0] Wgt_6_297, // sfix19_En18 
    input [18:0] Wgt_6_298, // sfix19_En18 
    input [18:0] Wgt_6_299, // sfix19_En18 
    input [18:0] Wgt_6_300, // sfix19_En18 
    input [18:0] Wgt_6_301, // sfix19_En18 
    input [18:0] Wgt_6_302, // sfix19_En18 
    input [18:0] Wgt_6_303, // sfix19_En18 
    input [18:0] Wgt_6_304, // sfix19_En18 
    input [18:0] Wgt_6_305, // sfix19_En18 
    input [18:0] Wgt_6_306, // sfix19_En18 
    input [18:0] Wgt_6_307, // sfix19_En18 
    input [18:0] Wgt_6_308, // sfix19_En18 
    input [18:0] Wgt_6_309, // sfix19_En18 
    input [18:0] Wgt_6_310, // sfix19_En18 
    input [18:0] Wgt_6_311, // sfix19_En18 
    input [18:0] Wgt_6_312, // sfix19_En18 
    input [18:0] Wgt_6_313, // sfix19_En18 
    input [18:0] Wgt_6_314, // sfix19_En18 
    input [18:0] Wgt_6_315, // sfix19_En18 
    input [18:0] Wgt_6_316, // sfix19_En18 
    input [18:0] Wgt_6_317, // sfix19_En18 
    input [18:0] Wgt_6_318, // sfix19_En18 
    input [18:0] Wgt_6_319, // sfix19_En18 
    input [18:0] Wgt_6_320, // sfix19_En18 
    input [18:0] Wgt_6_321, // sfix19_En18 
    input [18:0] Wgt_6_322, // sfix19_En18 
    input [18:0] Wgt_6_323, // sfix19_En18 
    input [18:0] Wgt_6_324, // sfix19_En18 
    input [18:0] Wgt_6_325, // sfix19_En18 
    input [18:0] Wgt_6_326, // sfix19_En18 
    input [18:0] Wgt_6_327, // sfix19_En18 
    input [18:0] Wgt_6_328, // sfix19_En18 
    input [18:0] Wgt_6_329, // sfix19_En18 
    input [18:0] Wgt_6_330, // sfix19_En18 
    input [18:0] Wgt_6_331, // sfix19_En18 
    input [18:0] Wgt_6_332, // sfix19_En18 
    input [18:0] Wgt_6_333, // sfix19_En18 
    input [18:0] Wgt_6_334, // sfix19_En18 
    input [18:0] Wgt_6_335, // sfix19_En18 
    input [18:0] Wgt_6_336, // sfix19_En18 
    input [18:0] Wgt_6_337, // sfix19_En18 
    input [18:0] Wgt_6_338, // sfix19_En18 
    input [18:0] Wgt_6_339, // sfix19_En18 
    input [18:0] Wgt_6_340, // sfix19_En18 
    input [18:0] Wgt_6_341, // sfix19_En18 
    input [18:0] Wgt_6_342, // sfix19_En18 
    input [18:0] Wgt_6_343, // sfix19_En18 
    input [18:0] Wgt_6_344, // sfix19_En18 
    input [18:0] Wgt_6_345, // sfix19_En18 
    input [18:0] Wgt_6_346, // sfix19_En18 
    input [18:0] Wgt_6_347, // sfix19_En18 
    input [18:0] Wgt_6_348, // sfix19_En18 
    input [18:0] Wgt_6_349, // sfix19_En18 
    input [18:0] Wgt_6_350, // sfix19_En18 
    input [18:0] Wgt_6_351, // sfix19_En18 
    input [18:0] Wgt_6_352, // sfix19_En18 
    input [18:0] Wgt_6_353, // sfix19_En18 
    input [18:0] Wgt_6_354, // sfix19_En18 
    input [18:0] Wgt_6_355, // sfix19_En18 
    input [18:0] Wgt_6_356, // sfix19_En18 
    input [18:0] Wgt_6_357, // sfix19_En18 
    input [18:0] Wgt_6_358, // sfix19_En18 
    input [18:0] Wgt_6_359, // sfix19_En18 
    input [18:0] Wgt_6_360, // sfix19_En18 
    input [18:0] Wgt_6_361, // sfix19_En18 
    input [18:0] Wgt_6_362, // sfix19_En18 
    input [18:0] Wgt_6_363, // sfix19_En18 
    input [18:0] Wgt_6_364, // sfix19_En18 
    input [18:0] Wgt_6_365, // sfix19_En18 
    input [18:0] Wgt_6_366, // sfix19_En18 
    input [18:0] Wgt_6_367, // sfix19_En18 
    input [18:0] Wgt_6_368, // sfix19_En18 
    input [18:0] Wgt_6_369, // sfix19_En18 
    input [18:0] Wgt_6_370, // sfix19_En18 
    input [18:0] Wgt_6_371, // sfix19_En18 
    input [18:0] Wgt_6_372, // sfix19_En18 
    input [18:0] Wgt_6_373, // sfix19_En18 
    input [18:0] Wgt_6_374, // sfix19_En18 
    input [18:0] Wgt_6_375, // sfix19_En18 
    input [18:0] Wgt_6_376, // sfix19_En18 
    input [18:0] Wgt_6_377, // sfix19_En18 
    input [18:0] Wgt_6_378, // sfix19_En18 
    input [18:0] Wgt_6_379, // sfix19_En18 
    input [18:0] Wgt_6_380, // sfix19_En18 
    input [18:0] Wgt_6_381, // sfix19_En18 
    input [18:0] Wgt_6_382, // sfix19_En18 
    input [18:0] Wgt_6_383, // sfix19_En18 
    input [18:0] Wgt_6_384, // sfix19_En18 
    input [18:0] Wgt_6_385, // sfix19_En18 
    input [18:0] Wgt_6_386, // sfix19_En18 
    input [18:0] Wgt_6_387, // sfix19_En18 
    input [18:0] Wgt_6_388, // sfix19_En18 
    input [18:0] Wgt_6_389, // sfix19_En18 
    input [18:0] Wgt_6_390, // sfix19_En18 
    input [18:0] Wgt_6_391, // sfix19_En18 
    input [18:0] Wgt_6_392, // sfix19_En18 
    input [18:0] Wgt_6_393, // sfix19_En18 
    input [18:0] Wgt_6_394, // sfix19_En18 
    input [18:0] Wgt_6_395, // sfix19_En18 
    input [18:0] Wgt_6_396, // sfix19_En18 
    input [18:0] Wgt_6_397, // sfix19_En18 
    input [18:0] Wgt_6_398, // sfix19_En18 
    input [18:0] Wgt_6_399, // sfix19_En18 
    input [18:0] Wgt_6_400, // sfix19_En18 
    input [18:0] Wgt_6_401, // sfix19_En18 
    input [18:0] Wgt_6_402, // sfix19_En18 
    input [18:0] Wgt_6_403, // sfix19_En18 
    input [18:0] Wgt_6_404, // sfix19_En18 
    input [18:0] Wgt_6_405, // sfix19_En18 
    input [18:0] Wgt_6_406, // sfix19_En18 
    input [18:0] Wgt_6_407, // sfix19_En18 
    input [18:0] Wgt_6_408, // sfix19_En18 
    input [18:0] Wgt_6_409, // sfix19_En18 
    input [18:0] Wgt_6_410, // sfix19_En18 
    input [18:0] Wgt_6_411, // sfix19_En18 
    input [18:0] Wgt_6_412, // sfix19_En18 
    input [18:0] Wgt_6_413, // sfix19_En18 
    input [18:0] Wgt_6_414, // sfix19_En18 
    input [18:0] Wgt_6_415, // sfix19_En18 
    input [18:0] Wgt_6_416, // sfix19_En18 
    input [18:0] Wgt_6_417, // sfix19_En18 
    input [18:0] Wgt_6_418, // sfix19_En18 
    input [18:0] Wgt_6_419, // sfix19_En18 
    input [18:0] Wgt_6_420, // sfix19_En18 
    input [18:0] Wgt_6_421, // sfix19_En18 
    input [18:0] Wgt_6_422, // sfix19_En18 
    input [18:0] Wgt_6_423, // sfix19_En18 
    input [18:0] Wgt_6_424, // sfix19_En18 
    input [18:0] Wgt_6_425, // sfix19_En18 
    input [18:0] Wgt_6_426, // sfix19_En18 
    input [18:0] Wgt_6_427, // sfix19_En18 
    input [18:0] Wgt_6_428, // sfix19_En18 
    input [18:0] Wgt_6_429, // sfix19_En18 
    input [18:0] Wgt_6_430, // sfix19_En18 
    input [18:0] Wgt_6_431, // sfix19_En18 
    input [18:0] Wgt_6_432, // sfix19_En18 
    input [18:0] Wgt_6_433, // sfix19_En18 
    input [18:0] Wgt_6_434, // sfix19_En18 
    input [18:0] Wgt_6_435, // sfix19_En18 
    input [18:0] Wgt_6_436, // sfix19_En18 
    input [18:0] Wgt_6_437, // sfix19_En18 
    input [18:0] Wgt_6_438, // sfix19_En18 
    input [18:0] Wgt_6_439, // sfix19_En18 
    input [18:0] Wgt_6_440, // sfix19_En18 
    input [18:0] Wgt_6_441, // sfix19_En18 
    input [18:0] Wgt_6_442, // sfix19_En18 
    input [18:0] Wgt_6_443, // sfix19_En18 
    input [18:0] Wgt_6_444, // sfix19_En18 
    input [18:0] Wgt_6_445, // sfix19_En18 
    input [18:0] Wgt_6_446, // sfix19_En18 
    input [18:0] Wgt_6_447, // sfix19_En18 
    input [18:0] Wgt_6_448, // sfix19_En18 
    input [18:0] Wgt_6_449, // sfix19_En18 
    input [18:0] Wgt_6_450, // sfix19_En18 
    input [18:0] Wgt_6_451, // sfix19_En18 
    input [18:0] Wgt_6_452, // sfix19_En18 
    input [18:0] Wgt_6_453, // sfix19_En18 
    input [18:0] Wgt_6_454, // sfix19_En18 
    input [18:0] Wgt_6_455, // sfix19_En18 
    input [18:0] Wgt_6_456, // sfix19_En18 
    input [18:0] Wgt_6_457, // sfix19_En18 
    input [18:0] Wgt_6_458, // sfix19_En18 
    input [18:0] Wgt_6_459, // sfix19_En18 
    input [18:0] Wgt_6_460, // sfix19_En18 
    input [18:0] Wgt_6_461, // sfix19_En18 
    input [18:0] Wgt_6_462, // sfix19_En18 
    input [18:0] Wgt_6_463, // sfix19_En18 
    input [18:0] Wgt_6_464, // sfix19_En18 
    input [18:0] Wgt_6_465, // sfix19_En18 
    input [18:0] Wgt_6_466, // sfix19_En18 
    input [18:0] Wgt_6_467, // sfix19_En18 
    input [18:0] Wgt_6_468, // sfix19_En18 
    input [18:0] Wgt_6_469, // sfix19_En18 
    input [18:0] Wgt_6_470, // sfix19_En18 
    input [18:0] Wgt_6_471, // sfix19_En18 
    input [18:0] Wgt_6_472, // sfix19_En18 
    input [18:0] Wgt_6_473, // sfix19_En18 
    input [18:0] Wgt_6_474, // sfix19_En18 
    input [18:0] Wgt_6_475, // sfix19_En18 
    input [18:0] Wgt_6_476, // sfix19_En18 
    input [18:0] Wgt_6_477, // sfix19_En18 
    input [18:0] Wgt_6_478, // sfix19_En18 
    input [18:0] Wgt_6_479, // sfix19_En18 
    input [18:0] Wgt_6_480, // sfix19_En18 
    input [18:0] Wgt_6_481, // sfix19_En18 
    input [18:0] Wgt_6_482, // sfix19_En18 
    input [18:0] Wgt_6_483, // sfix19_En18 
    input [18:0] Wgt_6_484, // sfix19_En18 
    input [18:0] Wgt_6_485, // sfix19_En18 
    input [18:0] Wgt_6_486, // sfix19_En18 
    input [18:0] Wgt_6_487, // sfix19_En18 
    input [18:0] Wgt_6_488, // sfix19_En18 
    input [18:0] Wgt_6_489, // sfix19_En18 
    input [18:0] Wgt_6_490, // sfix19_En18 
    input [18:0] Wgt_6_491, // sfix19_En18 
    input [18:0] Wgt_6_492, // sfix19_En18 
    input [18:0] Wgt_6_493, // sfix19_En18 
    input [18:0] Wgt_6_494, // sfix19_En18 
    input [18:0] Wgt_6_495, // sfix19_En18 
    input [18:0] Wgt_6_496, // sfix19_En18 
    input [18:0] Wgt_6_497, // sfix19_En18 
    input [18:0] Wgt_6_498, // sfix19_En18 
    input [18:0] Wgt_6_499, // sfix19_En18 
    input [18:0] Wgt_6_500, // sfix19_En18 
    input [18:0] Wgt_6_501, // sfix19_En18 
    input [18:0] Wgt_6_502, // sfix19_En18 
    input [18:0] Wgt_6_503, // sfix19_En18 
    input [18:0] Wgt_6_504, // sfix19_En18 
    input [18:0] Wgt_6_505, // sfix19_En18 
    input [18:0] Wgt_6_506, // sfix19_En18 
    input [18:0] Wgt_6_507, // sfix19_En18 
    input [18:0] Wgt_6_508, // sfix19_En18 
    input [18:0] Wgt_6_509, // sfix19_En18 
    input [18:0] Wgt_6_510, // sfix19_En18 
    input [18:0] Wgt_6_511, // sfix19_En18 
    input [18:0] Wgt_6_512, // sfix19_En18 
    input [18:0] Wgt_6_513, // sfix19_En18 
    input [18:0] Wgt_6_514, // sfix19_En18 
    input [18:0] Wgt_6_515, // sfix19_En18 
    input [18:0] Wgt_6_516, // sfix19_En18 
    input [18:0] Wgt_6_517, // sfix19_En18 
    input [18:0] Wgt_6_518, // sfix19_En18 
    input [18:0] Wgt_6_519, // sfix19_En18 
    input [18:0] Wgt_6_520, // sfix19_En18 
    input [18:0] Wgt_6_521, // sfix19_En18 
    input [18:0] Wgt_6_522, // sfix19_En18 
    input [18:0] Wgt_6_523, // sfix19_En18 
    input [18:0] Wgt_6_524, // sfix19_En18 
    input [18:0] Wgt_6_525, // sfix19_En18 
    input [18:0] Wgt_6_526, // sfix19_En18 
    input [18:0] Wgt_6_527, // sfix19_En18 
    input [18:0] Wgt_6_528, // sfix19_En18 
    input [18:0] Wgt_6_529, // sfix19_En18 
    input [18:0] Wgt_6_530, // sfix19_En18 
    input [18:0] Wgt_6_531, // sfix19_En18 
    input [18:0] Wgt_6_532, // sfix19_En18 
    input [18:0] Wgt_6_533, // sfix19_En18 
    input [18:0] Wgt_6_534, // sfix19_En18 
    input [18:0] Wgt_6_535, // sfix19_En18 
    input [18:0] Wgt_6_536, // sfix19_En18 
    input [18:0] Wgt_6_537, // sfix19_En18 
    input [18:0] Wgt_6_538, // sfix19_En18 
    input [18:0] Wgt_6_539, // sfix19_En18 
    input [18:0] Wgt_6_540, // sfix19_En18 
    input [18:0] Wgt_6_541, // sfix19_En18 
    input [18:0] Wgt_6_542, // sfix19_En18 
    input [18:0] Wgt_6_543, // sfix19_En18 
    input [18:0] Wgt_6_544, // sfix19_En18 
    input [18:0] Wgt_6_545, // sfix19_En18 
    input [18:0] Wgt_6_546, // sfix19_En18 
    input [18:0] Wgt_6_547, // sfix19_En18 
    input [18:0] Wgt_6_548, // sfix19_En18 
    input [18:0] Wgt_6_549, // sfix19_En18 
    input [18:0] Wgt_6_550, // sfix19_En18 
    input [18:0] Wgt_6_551, // sfix19_En18 
    input [18:0] Wgt_6_552, // sfix19_En18 
    input [18:0] Wgt_6_553, // sfix19_En18 
    input [18:0] Wgt_6_554, // sfix19_En18 
    input [18:0] Wgt_6_555, // sfix19_En18 
    input [18:0] Wgt_6_556, // sfix19_En18 
    input [18:0] Wgt_6_557, // sfix19_En18 
    input [18:0] Wgt_6_558, // sfix19_En18 
    input [18:0] Wgt_6_559, // sfix19_En18 
    input [18:0] Wgt_6_560, // sfix19_En18 
    input [18:0] Wgt_6_561, // sfix19_En18 
    input [18:0] Wgt_6_562, // sfix19_En18 
    input [18:0] Wgt_6_563, // sfix19_En18 
    input [18:0] Wgt_6_564, // sfix19_En18 
    input [18:0] Wgt_6_565, // sfix19_En18 
    input [18:0] Wgt_6_566, // sfix19_En18 
    input [18:0] Wgt_6_567, // sfix19_En18 
    input [18:0] Wgt_6_568, // sfix19_En18 
    input [18:0] Wgt_6_569, // sfix19_En18 
    input [18:0] Wgt_6_570, // sfix19_En18 
    input [18:0] Wgt_6_571, // sfix19_En18 
    input [18:0] Wgt_6_572, // sfix19_En18 
    input [18:0] Wgt_6_573, // sfix19_En18 
    input [18:0] Wgt_6_574, // sfix19_En18 
    input [18:0] Wgt_6_575, // sfix19_En18 
    input [18:0] Wgt_6_576, // sfix19_En18 
    input [18:0] Wgt_6_577, // sfix19_En18 
    input [18:0] Wgt_6_578, // sfix19_En18 
    input [18:0] Wgt_6_579, // sfix19_En18 
    input [18:0] Wgt_6_580, // sfix19_En18 
    input [18:0] Wgt_6_581, // sfix19_En18 
    input [18:0] Wgt_6_582, // sfix19_En18 
    input [18:0] Wgt_6_583, // sfix19_En18 
    input [18:0] Wgt_6_584, // sfix19_En18 
    input [18:0] Wgt_6_585, // sfix19_En18 
    input [18:0] Wgt_6_586, // sfix19_En18 
    input [18:0] Wgt_6_587, // sfix19_En18 
    input [18:0] Wgt_6_588, // sfix19_En18 
    input [18:0] Wgt_6_589, // sfix19_En18 
    input [18:0] Wgt_6_590, // sfix19_En18 
    input [18:0] Wgt_6_591, // sfix19_En18 
    input [18:0] Wgt_6_592, // sfix19_En18 
    input [18:0] Wgt_6_593, // sfix19_En18 
    input [18:0] Wgt_6_594, // sfix19_En18 
    input [18:0] Wgt_6_595, // sfix19_En18 
    input [18:0] Wgt_6_596, // sfix19_En18 
    input [18:0] Wgt_6_597, // sfix19_En18 
    input [18:0] Wgt_6_598, // sfix19_En18 
    input [18:0] Wgt_6_599, // sfix19_En18 
    input [18:0] Wgt_6_600, // sfix19_En18 
    input [18:0] Wgt_6_601, // sfix19_En18 
    input [18:0] Wgt_6_602, // sfix19_En18 
    input [18:0] Wgt_6_603, // sfix19_En18 
    input [18:0] Wgt_6_604, // sfix19_En18 
    input [18:0] Wgt_6_605, // sfix19_En18 
    input [18:0] Wgt_6_606, // sfix19_En18 
    input [18:0] Wgt_6_607, // sfix19_En18 
    input [18:0] Wgt_6_608, // sfix19_En18 
    input [18:0] Wgt_6_609, // sfix19_En18 
    input [18:0] Wgt_6_610, // sfix19_En18 
    input [18:0] Wgt_6_611, // sfix19_En18 
    input [18:0] Wgt_6_612, // sfix19_En18 
    input [18:0] Wgt_6_613, // sfix19_En18 
    input [18:0] Wgt_6_614, // sfix19_En18 
    input [18:0] Wgt_6_615, // sfix19_En18 
    input [18:0] Wgt_6_616, // sfix19_En18 
    input [18:0] Wgt_6_617, // sfix19_En18 
    input [18:0] Wgt_6_618, // sfix19_En18 
    input [18:0] Wgt_6_619, // sfix19_En18 
    input [18:0] Wgt_6_620, // sfix19_En18 
    input [18:0] Wgt_6_621, // sfix19_En18 
    input [18:0] Wgt_6_622, // sfix19_En18 
    input [18:0] Wgt_6_623, // sfix19_En18 
    input [18:0] Wgt_6_624, // sfix19_En18 
    input [18:0] Wgt_6_625, // sfix19_En18 
    input [18:0] Wgt_6_626, // sfix19_En18 
    input [18:0] Wgt_6_627, // sfix19_En18 
    input [18:0] Wgt_6_628, // sfix19_En18 
    input [18:0] Wgt_6_629, // sfix19_En18 
    input [18:0] Wgt_6_630, // sfix19_En18 
    input [18:0] Wgt_6_631, // sfix19_En18 
    input [18:0] Wgt_6_632, // sfix19_En18 
    input [18:0] Wgt_6_633, // sfix19_En18 
    input [18:0] Wgt_6_634, // sfix19_En18 
    input [18:0] Wgt_6_635, // sfix19_En18 
    input [18:0] Wgt_6_636, // sfix19_En18 
    input [18:0] Wgt_6_637, // sfix19_En18 
    input [18:0] Wgt_6_638, // sfix19_En18 
    input [18:0] Wgt_6_639, // sfix19_En18 
    input [18:0] Wgt_6_640, // sfix19_En18 
    input [18:0] Wgt_6_641, // sfix19_En18 
    input [18:0] Wgt_6_642, // sfix19_En18 
    input [18:0] Wgt_6_643, // sfix19_En18 
    input [18:0] Wgt_6_644, // sfix19_En18 
    input [18:0] Wgt_6_645, // sfix19_En18 
    input [18:0] Wgt_6_646, // sfix19_En18 
    input [18:0] Wgt_6_647, // sfix19_En18 
    input [18:0] Wgt_6_648, // sfix19_En18 
    input [18:0] Wgt_6_649, // sfix19_En18 
    input [18:0] Wgt_6_650, // sfix19_En18 
    input [18:0] Wgt_6_651, // sfix19_En18 
    input [18:0] Wgt_6_652, // sfix19_En18 
    input [18:0] Wgt_6_653, // sfix19_En18 
    input [18:0] Wgt_6_654, // sfix19_En18 
    input [18:0] Wgt_6_655, // sfix19_En18 
    input [18:0] Wgt_6_656, // sfix19_En18 
    input [18:0] Wgt_6_657, // sfix19_En18 
    input [18:0] Wgt_6_658, // sfix19_En18 
    input [18:0] Wgt_6_659, // sfix19_En18 
    input [18:0] Wgt_6_660, // sfix19_En18 
    input [18:0] Wgt_6_661, // sfix19_En18 
    input [18:0] Wgt_6_662, // sfix19_En18 
    input [18:0] Wgt_6_663, // sfix19_En18 
    input [18:0] Wgt_6_664, // sfix19_En18 
    input [18:0] Wgt_6_665, // sfix19_En18 
    input [18:0] Wgt_6_666, // sfix19_En18 
    input [18:0] Wgt_6_667, // sfix19_En18 
    input [18:0] Wgt_6_668, // sfix19_En18 
    input [18:0] Wgt_6_669, // sfix19_En18 
    input [18:0] Wgt_6_670, // sfix19_En18 
    input [18:0] Wgt_6_671, // sfix19_En18 
    input [18:0] Wgt_6_672, // sfix19_En18 
    input [18:0] Wgt_6_673, // sfix19_En18 
    input [18:0] Wgt_6_674, // sfix19_En18 
    input [18:0] Wgt_6_675, // sfix19_En18 
    input [18:0] Wgt_6_676, // sfix19_En18 
    input [18:0] Wgt_6_677, // sfix19_En18 
    input [18:0] Wgt_6_678, // sfix19_En18 
    input [18:0] Wgt_6_679, // sfix19_En18 
    input [18:0] Wgt_6_680, // sfix19_En18 
    input [18:0] Wgt_6_681, // sfix19_En18 
    input [18:0] Wgt_6_682, // sfix19_En18 
    input [18:0] Wgt_6_683, // sfix19_En18 
    input [18:0] Wgt_6_684, // sfix19_En18 
    input [18:0] Wgt_6_685, // sfix19_En18 
    input [18:0] Wgt_6_686, // sfix19_En18 
    input [18:0] Wgt_6_687, // sfix19_En18 
    input [18:0] Wgt_6_688, // sfix19_En18 
    input [18:0] Wgt_6_689, // sfix19_En18 
    input [18:0] Wgt_6_690, // sfix19_En18 
    input [18:0] Wgt_6_691, // sfix19_En18 
    input [18:0] Wgt_6_692, // sfix19_En18 
    input [18:0] Wgt_6_693, // sfix19_En18 
    input [18:0] Wgt_6_694, // sfix19_En18 
    input [18:0] Wgt_6_695, // sfix19_En18 
    input [18:0] Wgt_6_696, // sfix19_En18 
    input [18:0] Wgt_6_697, // sfix19_En18 
    input [18:0] Wgt_6_698, // sfix19_En18 
    input [18:0] Wgt_6_699, // sfix19_En18 
    input [18:0] Wgt_6_700, // sfix19_En18 
    input [18:0] Wgt_6_701, // sfix19_En18 
    input [18:0] Wgt_6_702, // sfix19_En18 
    input [18:0] Wgt_6_703, // sfix19_En18 
    input [18:0] Wgt_6_704, // sfix19_En18 
    input [18:0] Wgt_6_705, // sfix19_En18 
    input [18:0] Wgt_6_706, // sfix19_En18 
    input [18:0] Wgt_6_707, // sfix19_En18 
    input [18:0] Wgt_6_708, // sfix19_En18 
    input [18:0] Wgt_6_709, // sfix19_En18 
    input [18:0] Wgt_6_710, // sfix19_En18 
    input [18:0] Wgt_6_711, // sfix19_En18 
    input [18:0] Wgt_6_712, // sfix19_En18 
    input [18:0] Wgt_6_713, // sfix19_En18 
    input [18:0] Wgt_6_714, // sfix19_En18 
    input [18:0] Wgt_6_715, // sfix19_En18 
    input [18:0] Wgt_6_716, // sfix19_En18 
    input [18:0] Wgt_6_717, // sfix19_En18 
    input [18:0] Wgt_6_718, // sfix19_En18 
    input [18:0] Wgt_6_719, // sfix19_En18 
    input [18:0] Wgt_6_720, // sfix19_En18 
    input [18:0] Wgt_6_721, // sfix19_En18 
    input [18:0] Wgt_6_722, // sfix19_En18 
    input [18:0] Wgt_6_723, // sfix19_En18 
    input [18:0] Wgt_6_724, // sfix19_En18 
    input [18:0] Wgt_6_725, // sfix19_En18 
    input [18:0] Wgt_6_726, // sfix19_En18 
    input [18:0] Wgt_6_727, // sfix19_En18 
    input [18:0] Wgt_6_728, // sfix19_En18 
    input [18:0] Wgt_6_729, // sfix19_En18 
    input [18:0] Wgt_6_730, // sfix19_En18 
    input [18:0] Wgt_6_731, // sfix19_En18 
    input [18:0] Wgt_6_732, // sfix19_En18 
    input [18:0] Wgt_6_733, // sfix19_En18 
    input [18:0] Wgt_6_734, // sfix19_En18 
    input [18:0] Wgt_6_735, // sfix19_En18 
    input [18:0] Wgt_6_736, // sfix19_En18 
    input [18:0] Wgt_6_737, // sfix19_En18 
    input [18:0] Wgt_6_738, // sfix19_En18 
    input [18:0] Wgt_6_739, // sfix19_En18 
    input [18:0] Wgt_6_740, // sfix19_En18 
    input [18:0] Wgt_6_741, // sfix19_En18 
    input [18:0] Wgt_6_742, // sfix19_En18 
    input [18:0] Wgt_6_743, // sfix19_En18 
    input [18:0] Wgt_6_744, // sfix19_En18 
    input [18:0] Wgt_6_745, // sfix19_En18 
    input [18:0] Wgt_6_746, // sfix19_En18 
    input [18:0] Wgt_6_747, // sfix19_En18 
    input [18:0] Wgt_6_748, // sfix19_En18 
    input [18:0] Wgt_6_749, // sfix19_En18 
    input [18:0] Wgt_6_750, // sfix19_En18 
    input [18:0] Wgt_6_751, // sfix19_En18 
    input [18:0] Wgt_6_752, // sfix19_En18 
    input [18:0] Wgt_6_753, // sfix19_En18 
    input [18:0] Wgt_6_754, // sfix19_En18 
    input [18:0] Wgt_6_755, // sfix19_En18 
    input [18:0] Wgt_6_756, // sfix19_En18 
    input [18:0] Wgt_6_757, // sfix19_En18 
    input [18:0] Wgt_6_758, // sfix19_En18 
    input [18:0] Wgt_6_759, // sfix19_En18 
    input [18:0] Wgt_6_760, // sfix19_En18 
    input [18:0] Wgt_6_761, // sfix19_En18 
    input [18:0] Wgt_6_762, // sfix19_En18 
    input [18:0] Wgt_6_763, // sfix19_En18 
    input [18:0] Wgt_6_764, // sfix19_En18 
    input [18:0] Wgt_6_765, // sfix19_En18 
    input [18:0] Wgt_6_766, // sfix19_En18 
    input [18:0] Wgt_6_767, // sfix19_En18 
    input [18:0] Wgt_6_768, // sfix19_En18 
    input [18:0] Wgt_6_769, // sfix19_En18 
    input [18:0] Wgt_6_770, // sfix19_En18 
    input [18:0] Wgt_6_771, // sfix19_En18 
    input [18:0] Wgt_6_772, // sfix19_En18 
    input [18:0] Wgt_6_773, // sfix19_En18 
    input [18:0] Wgt_6_774, // sfix19_En18 
    input [18:0] Wgt_6_775, // sfix19_En18 
    input [18:0] Wgt_6_776, // sfix19_En18 
    input [18:0] Wgt_6_777, // sfix19_En18 
    input [18:0] Wgt_6_778, // sfix19_En18 
    input [18:0] Wgt_6_779, // sfix19_En18 
    input [18:0] Wgt_6_780, // sfix19_En18 
    input [18:0] Wgt_6_781, // sfix19_En18 
    input [18:0] Wgt_6_782, // sfix19_En18 
    input [18:0] Wgt_6_783, // sfix19_En18 
    input [18:0] Wgt_6_784, // sfix19_En18 
    input [18:0] Wgt_7_0, // sfix19_En18 
    input [18:0] Wgt_7_1, // sfix19_En18 
    input [18:0] Wgt_7_2, // sfix19_En18 
    input [18:0] Wgt_7_3, // sfix19_En18 
    input [18:0] Wgt_7_4, // sfix19_En18 
    input [18:0] Wgt_7_5, // sfix19_En18 
    input [18:0] Wgt_7_6, // sfix19_En18 
    input [18:0] Wgt_7_7, // sfix19_En18 
    input [18:0] Wgt_7_8, // sfix19_En18 
    input [18:0] Wgt_7_9, // sfix19_En18 
    input [18:0] Wgt_7_10, // sfix19_En18 
    input [18:0] Wgt_7_11, // sfix19_En18 
    input [18:0] Wgt_7_12, // sfix19_En18 
    input [18:0] Wgt_7_13, // sfix19_En18 
    input [18:0] Wgt_7_14, // sfix19_En18 
    input [18:0] Wgt_7_15, // sfix19_En18 
    input [18:0] Wgt_7_16, // sfix19_En18 
    input [18:0] Wgt_7_17, // sfix19_En18 
    input [18:0] Wgt_7_18, // sfix19_En18 
    input [18:0] Wgt_7_19, // sfix19_En18 
    input [18:0] Wgt_7_20, // sfix19_En18 
    input [18:0] Wgt_7_21, // sfix19_En18 
    input [18:0] Wgt_7_22, // sfix19_En18 
    input [18:0] Wgt_7_23, // sfix19_En18 
    input [18:0] Wgt_7_24, // sfix19_En18 
    input [18:0] Wgt_7_25, // sfix19_En18 
    input [18:0] Wgt_7_26, // sfix19_En18 
    input [18:0] Wgt_7_27, // sfix19_En18 
    input [18:0] Wgt_7_28, // sfix19_En18 
    input [18:0] Wgt_7_29, // sfix19_En18 
    input [18:0] Wgt_7_30, // sfix19_En18 
    input [18:0] Wgt_7_31, // sfix19_En18 
    input [18:0] Wgt_7_32, // sfix19_En18 
    input [18:0] Wgt_7_33, // sfix19_En18 
    input [18:0] Wgt_7_34, // sfix19_En18 
    input [18:0] Wgt_7_35, // sfix19_En18 
    input [18:0] Wgt_7_36, // sfix19_En18 
    input [18:0] Wgt_7_37, // sfix19_En18 
    input [18:0] Wgt_7_38, // sfix19_En18 
    input [18:0] Wgt_7_39, // sfix19_En18 
    input [18:0] Wgt_7_40, // sfix19_En18 
    input [18:0] Wgt_7_41, // sfix19_En18 
    input [18:0] Wgt_7_42, // sfix19_En18 
    input [18:0] Wgt_7_43, // sfix19_En18 
    input [18:0] Wgt_7_44, // sfix19_En18 
    input [18:0] Wgt_7_45, // sfix19_En18 
    input [18:0] Wgt_7_46, // sfix19_En18 
    input [18:0] Wgt_7_47, // sfix19_En18 
    input [18:0] Wgt_7_48, // sfix19_En18 
    input [18:0] Wgt_7_49, // sfix19_En18 
    input [18:0] Wgt_7_50, // sfix19_En18 
    input [18:0] Wgt_7_51, // sfix19_En18 
    input [18:0] Wgt_7_52, // sfix19_En18 
    input [18:0] Wgt_7_53, // sfix19_En18 
    input [18:0] Wgt_7_54, // sfix19_En18 
    input [18:0] Wgt_7_55, // sfix19_En18 
    input [18:0] Wgt_7_56, // sfix19_En18 
    input [18:0] Wgt_7_57, // sfix19_En18 
    input [18:0] Wgt_7_58, // sfix19_En18 
    input [18:0] Wgt_7_59, // sfix19_En18 
    input [18:0] Wgt_7_60, // sfix19_En18 
    input [18:0] Wgt_7_61, // sfix19_En18 
    input [18:0] Wgt_7_62, // sfix19_En18 
    input [18:0] Wgt_7_63, // sfix19_En18 
    input [18:0] Wgt_7_64, // sfix19_En18 
    input [18:0] Wgt_7_65, // sfix19_En18 
    input [18:0] Wgt_7_66, // sfix19_En18 
    input [18:0] Wgt_7_67, // sfix19_En18 
    input [18:0] Wgt_7_68, // sfix19_En18 
    input [18:0] Wgt_7_69, // sfix19_En18 
    input [18:0] Wgt_7_70, // sfix19_En18 
    input [18:0] Wgt_7_71, // sfix19_En18 
    input [18:0] Wgt_7_72, // sfix19_En18 
    input [18:0] Wgt_7_73, // sfix19_En18 
    input [18:0] Wgt_7_74, // sfix19_En18 
    input [18:0] Wgt_7_75, // sfix19_En18 
    input [18:0] Wgt_7_76, // sfix19_En18 
    input [18:0] Wgt_7_77, // sfix19_En18 
    input [18:0] Wgt_7_78, // sfix19_En18 
    input [18:0] Wgt_7_79, // sfix19_En18 
    input [18:0] Wgt_7_80, // sfix19_En18 
    input [18:0] Wgt_7_81, // sfix19_En18 
    input [18:0] Wgt_7_82, // sfix19_En18 
    input [18:0] Wgt_7_83, // sfix19_En18 
    input [18:0] Wgt_7_84, // sfix19_En18 
    input [18:0] Wgt_7_85, // sfix19_En18 
    input [18:0] Wgt_7_86, // sfix19_En18 
    input [18:0] Wgt_7_87, // sfix19_En18 
    input [18:0] Wgt_7_88, // sfix19_En18 
    input [18:0] Wgt_7_89, // sfix19_En18 
    input [18:0] Wgt_7_90, // sfix19_En18 
    input [18:0] Wgt_7_91, // sfix19_En18 
    input [18:0] Wgt_7_92, // sfix19_En18 
    input [18:0] Wgt_7_93, // sfix19_En18 
    input [18:0] Wgt_7_94, // sfix19_En18 
    input [18:0] Wgt_7_95, // sfix19_En18 
    input [18:0] Wgt_7_96, // sfix19_En18 
    input [18:0] Wgt_7_97, // sfix19_En18 
    input [18:0] Wgt_7_98, // sfix19_En18 
    input [18:0] Wgt_7_99, // sfix19_En18 
    input [18:0] Wgt_7_100, // sfix19_En18 
    input [18:0] Wgt_7_101, // sfix19_En18 
    input [18:0] Wgt_7_102, // sfix19_En18 
    input [18:0] Wgt_7_103, // sfix19_En18 
    input [18:0] Wgt_7_104, // sfix19_En18 
    input [18:0] Wgt_7_105, // sfix19_En18 
    input [18:0] Wgt_7_106, // sfix19_En18 
    input [18:0] Wgt_7_107, // sfix19_En18 
    input [18:0] Wgt_7_108, // sfix19_En18 
    input [18:0] Wgt_7_109, // sfix19_En18 
    input [18:0] Wgt_7_110, // sfix19_En18 
    input [18:0] Wgt_7_111, // sfix19_En18 
    input [18:0] Wgt_7_112, // sfix19_En18 
    input [18:0] Wgt_7_113, // sfix19_En18 
    input [18:0] Wgt_7_114, // sfix19_En18 
    input [18:0] Wgt_7_115, // sfix19_En18 
    input [18:0] Wgt_7_116, // sfix19_En18 
    input [18:0] Wgt_7_117, // sfix19_En18 
    input [18:0] Wgt_7_118, // sfix19_En18 
    input [18:0] Wgt_7_119, // sfix19_En18 
    input [18:0] Wgt_7_120, // sfix19_En18 
    input [18:0] Wgt_7_121, // sfix19_En18 
    input [18:0] Wgt_7_122, // sfix19_En18 
    input [18:0] Wgt_7_123, // sfix19_En18 
    input [18:0] Wgt_7_124, // sfix19_En18 
    input [18:0] Wgt_7_125, // sfix19_En18 
    input [18:0] Wgt_7_126, // sfix19_En18 
    input [18:0] Wgt_7_127, // sfix19_En18 
    input [18:0] Wgt_7_128, // sfix19_En18 
    input [18:0] Wgt_7_129, // sfix19_En18 
    input [18:0] Wgt_7_130, // sfix19_En18 
    input [18:0] Wgt_7_131, // sfix19_En18 
    input [18:0] Wgt_7_132, // sfix19_En18 
    input [18:0] Wgt_7_133, // sfix19_En18 
    input [18:0] Wgt_7_134, // sfix19_En18 
    input [18:0] Wgt_7_135, // sfix19_En18 
    input [18:0] Wgt_7_136, // sfix19_En18 
    input [18:0] Wgt_7_137, // sfix19_En18 
    input [18:0] Wgt_7_138, // sfix19_En18 
    input [18:0] Wgt_7_139, // sfix19_En18 
    input [18:0] Wgt_7_140, // sfix19_En18 
    input [18:0] Wgt_7_141, // sfix19_En18 
    input [18:0] Wgt_7_142, // sfix19_En18 
    input [18:0] Wgt_7_143, // sfix19_En18 
    input [18:0] Wgt_7_144, // sfix19_En18 
    input [18:0] Wgt_7_145, // sfix19_En18 
    input [18:0] Wgt_7_146, // sfix19_En18 
    input [18:0] Wgt_7_147, // sfix19_En18 
    input [18:0] Wgt_7_148, // sfix19_En18 
    input [18:0] Wgt_7_149, // sfix19_En18 
    input [18:0] Wgt_7_150, // sfix19_En18 
    input [18:0] Wgt_7_151, // sfix19_En18 
    input [18:0] Wgt_7_152, // sfix19_En18 
    input [18:0] Wgt_7_153, // sfix19_En18 
    input [18:0] Wgt_7_154, // sfix19_En18 
    input [18:0] Wgt_7_155, // sfix19_En18 
    input [18:0] Wgt_7_156, // sfix19_En18 
    input [18:0] Wgt_7_157, // sfix19_En18 
    input [18:0] Wgt_7_158, // sfix19_En18 
    input [18:0] Wgt_7_159, // sfix19_En18 
    input [18:0] Wgt_7_160, // sfix19_En18 
    input [18:0] Wgt_7_161, // sfix19_En18 
    input [18:0] Wgt_7_162, // sfix19_En18 
    input [18:0] Wgt_7_163, // sfix19_En18 
    input [18:0] Wgt_7_164, // sfix19_En18 
    input [18:0] Wgt_7_165, // sfix19_En18 
    input [18:0] Wgt_7_166, // sfix19_En18 
    input [18:0] Wgt_7_167, // sfix19_En18 
    input [18:0] Wgt_7_168, // sfix19_En18 
    input [18:0] Wgt_7_169, // sfix19_En18 
    input [18:0] Wgt_7_170, // sfix19_En18 
    input [18:0] Wgt_7_171, // sfix19_En18 
    input [18:0] Wgt_7_172, // sfix19_En18 
    input [18:0] Wgt_7_173, // sfix19_En18 
    input [18:0] Wgt_7_174, // sfix19_En18 
    input [18:0] Wgt_7_175, // sfix19_En18 
    input [18:0] Wgt_7_176, // sfix19_En18 
    input [18:0] Wgt_7_177, // sfix19_En18 
    input [18:0] Wgt_7_178, // sfix19_En18 
    input [18:0] Wgt_7_179, // sfix19_En18 
    input [18:0] Wgt_7_180, // sfix19_En18 
    input [18:0] Wgt_7_181, // sfix19_En18 
    input [18:0] Wgt_7_182, // sfix19_En18 
    input [18:0] Wgt_7_183, // sfix19_En18 
    input [18:0] Wgt_7_184, // sfix19_En18 
    input [18:0] Wgt_7_185, // sfix19_En18 
    input [18:0] Wgt_7_186, // sfix19_En18 
    input [18:0] Wgt_7_187, // sfix19_En18 
    input [18:0] Wgt_7_188, // sfix19_En18 
    input [18:0] Wgt_7_189, // sfix19_En18 
    input [18:0] Wgt_7_190, // sfix19_En18 
    input [18:0] Wgt_7_191, // sfix19_En18 
    input [18:0] Wgt_7_192, // sfix19_En18 
    input [18:0] Wgt_7_193, // sfix19_En18 
    input [18:0] Wgt_7_194, // sfix19_En18 
    input [18:0] Wgt_7_195, // sfix19_En18 
    input [18:0] Wgt_7_196, // sfix19_En18 
    input [18:0] Wgt_7_197, // sfix19_En18 
    input [18:0] Wgt_7_198, // sfix19_En18 
    input [18:0] Wgt_7_199, // sfix19_En18 
    input [18:0] Wgt_7_200, // sfix19_En18 
    input [18:0] Wgt_7_201, // sfix19_En18 
    input [18:0] Wgt_7_202, // sfix19_En18 
    input [18:0] Wgt_7_203, // sfix19_En18 
    input [18:0] Wgt_7_204, // sfix19_En18 
    input [18:0] Wgt_7_205, // sfix19_En18 
    input [18:0] Wgt_7_206, // sfix19_En18 
    input [18:0] Wgt_7_207, // sfix19_En18 
    input [18:0] Wgt_7_208, // sfix19_En18 
    input [18:0] Wgt_7_209, // sfix19_En18 
    input [18:0] Wgt_7_210, // sfix19_En18 
    input [18:0] Wgt_7_211, // sfix19_En18 
    input [18:0] Wgt_7_212, // sfix19_En18 
    input [18:0] Wgt_7_213, // sfix19_En18 
    input [18:0] Wgt_7_214, // sfix19_En18 
    input [18:0] Wgt_7_215, // sfix19_En18 
    input [18:0] Wgt_7_216, // sfix19_En18 
    input [18:0] Wgt_7_217, // sfix19_En18 
    input [18:0] Wgt_7_218, // sfix19_En18 
    input [18:0] Wgt_7_219, // sfix19_En18 
    input [18:0] Wgt_7_220, // sfix19_En18 
    input [18:0] Wgt_7_221, // sfix19_En18 
    input [18:0] Wgt_7_222, // sfix19_En18 
    input [18:0] Wgt_7_223, // sfix19_En18 
    input [18:0] Wgt_7_224, // sfix19_En18 
    input [18:0] Wgt_7_225, // sfix19_En18 
    input [18:0] Wgt_7_226, // sfix19_En18 
    input [18:0] Wgt_7_227, // sfix19_En18 
    input [18:0] Wgt_7_228, // sfix19_En18 
    input [18:0] Wgt_7_229, // sfix19_En18 
    input [18:0] Wgt_7_230, // sfix19_En18 
    input [18:0] Wgt_7_231, // sfix19_En18 
    input [18:0] Wgt_7_232, // sfix19_En18 
    input [18:0] Wgt_7_233, // sfix19_En18 
    input [18:0] Wgt_7_234, // sfix19_En18 
    input [18:0] Wgt_7_235, // sfix19_En18 
    input [18:0] Wgt_7_236, // sfix19_En18 
    input [18:0] Wgt_7_237, // sfix19_En18 
    input [18:0] Wgt_7_238, // sfix19_En18 
    input [18:0] Wgt_7_239, // sfix19_En18 
    input [18:0] Wgt_7_240, // sfix19_En18 
    input [18:0] Wgt_7_241, // sfix19_En18 
    input [18:0] Wgt_7_242, // sfix19_En18 
    input [18:0] Wgt_7_243, // sfix19_En18 
    input [18:0] Wgt_7_244, // sfix19_En18 
    input [18:0] Wgt_7_245, // sfix19_En18 
    input [18:0] Wgt_7_246, // sfix19_En18 
    input [18:0] Wgt_7_247, // sfix19_En18 
    input [18:0] Wgt_7_248, // sfix19_En18 
    input [18:0] Wgt_7_249, // sfix19_En18 
    input [18:0] Wgt_7_250, // sfix19_En18 
    input [18:0] Wgt_7_251, // sfix19_En18 
    input [18:0] Wgt_7_252, // sfix19_En18 
    input [18:0] Wgt_7_253, // sfix19_En18 
    input [18:0] Wgt_7_254, // sfix19_En18 
    input [18:0] Wgt_7_255, // sfix19_En18 
    input [18:0] Wgt_7_256, // sfix19_En18 
    input [18:0] Wgt_7_257, // sfix19_En18 
    input [18:0] Wgt_7_258, // sfix19_En18 
    input [18:0] Wgt_7_259, // sfix19_En18 
    input [18:0] Wgt_7_260, // sfix19_En18 
    input [18:0] Wgt_7_261, // sfix19_En18 
    input [18:0] Wgt_7_262, // sfix19_En18 
    input [18:0] Wgt_7_263, // sfix19_En18 
    input [18:0] Wgt_7_264, // sfix19_En18 
    input [18:0] Wgt_7_265, // sfix19_En18 
    input [18:0] Wgt_7_266, // sfix19_En18 
    input [18:0] Wgt_7_267, // sfix19_En18 
    input [18:0] Wgt_7_268, // sfix19_En18 
    input [18:0] Wgt_7_269, // sfix19_En18 
    input [18:0] Wgt_7_270, // sfix19_En18 
    input [18:0] Wgt_7_271, // sfix19_En18 
    input [18:0] Wgt_7_272, // sfix19_En18 
    input [18:0] Wgt_7_273, // sfix19_En18 
    input [18:0] Wgt_7_274, // sfix19_En18 
    input [18:0] Wgt_7_275, // sfix19_En18 
    input [18:0] Wgt_7_276, // sfix19_En18 
    input [18:0] Wgt_7_277, // sfix19_En18 
    input [18:0] Wgt_7_278, // sfix19_En18 
    input [18:0] Wgt_7_279, // sfix19_En18 
    input [18:0] Wgt_7_280, // sfix19_En18 
    input [18:0] Wgt_7_281, // sfix19_En18 
    input [18:0] Wgt_7_282, // sfix19_En18 
    input [18:0] Wgt_7_283, // sfix19_En18 
    input [18:0] Wgt_7_284, // sfix19_En18 
    input [18:0] Wgt_7_285, // sfix19_En18 
    input [18:0] Wgt_7_286, // sfix19_En18 
    input [18:0] Wgt_7_287, // sfix19_En18 
    input [18:0] Wgt_7_288, // sfix19_En18 
    input [18:0] Wgt_7_289, // sfix19_En18 
    input [18:0] Wgt_7_290, // sfix19_En18 
    input [18:0] Wgt_7_291, // sfix19_En18 
    input [18:0] Wgt_7_292, // sfix19_En18 
    input [18:0] Wgt_7_293, // sfix19_En18 
    input [18:0] Wgt_7_294, // sfix19_En18 
    input [18:0] Wgt_7_295, // sfix19_En18 
    input [18:0] Wgt_7_296, // sfix19_En18 
    input [18:0] Wgt_7_297, // sfix19_En18 
    input [18:0] Wgt_7_298, // sfix19_En18 
    input [18:0] Wgt_7_299, // sfix19_En18 
    input [18:0] Wgt_7_300, // sfix19_En18 
    input [18:0] Wgt_7_301, // sfix19_En18 
    input [18:0] Wgt_7_302, // sfix19_En18 
    input [18:0] Wgt_7_303, // sfix19_En18 
    input [18:0] Wgt_7_304, // sfix19_En18 
    input [18:0] Wgt_7_305, // sfix19_En18 
    input [18:0] Wgt_7_306, // sfix19_En18 
    input [18:0] Wgt_7_307, // sfix19_En18 
    input [18:0] Wgt_7_308, // sfix19_En18 
    input [18:0] Wgt_7_309, // sfix19_En18 
    input [18:0] Wgt_7_310, // sfix19_En18 
    input [18:0] Wgt_7_311, // sfix19_En18 
    input [18:0] Wgt_7_312, // sfix19_En18 
    input [18:0] Wgt_7_313, // sfix19_En18 
    input [18:0] Wgt_7_314, // sfix19_En18 
    input [18:0] Wgt_7_315, // sfix19_En18 
    input [18:0] Wgt_7_316, // sfix19_En18 
    input [18:0] Wgt_7_317, // sfix19_En18 
    input [18:0] Wgt_7_318, // sfix19_En18 
    input [18:0] Wgt_7_319, // sfix19_En18 
    input [18:0] Wgt_7_320, // sfix19_En18 
    input [18:0] Wgt_7_321, // sfix19_En18 
    input [18:0] Wgt_7_322, // sfix19_En18 
    input [18:0] Wgt_7_323, // sfix19_En18 
    input [18:0] Wgt_7_324, // sfix19_En18 
    input [18:0] Wgt_7_325, // sfix19_En18 
    input [18:0] Wgt_7_326, // sfix19_En18 
    input [18:0] Wgt_7_327, // sfix19_En18 
    input [18:0] Wgt_7_328, // sfix19_En18 
    input [18:0] Wgt_7_329, // sfix19_En18 
    input [18:0] Wgt_7_330, // sfix19_En18 
    input [18:0] Wgt_7_331, // sfix19_En18 
    input [18:0] Wgt_7_332, // sfix19_En18 
    input [18:0] Wgt_7_333, // sfix19_En18 
    input [18:0] Wgt_7_334, // sfix19_En18 
    input [18:0] Wgt_7_335, // sfix19_En18 
    input [18:0] Wgt_7_336, // sfix19_En18 
    input [18:0] Wgt_7_337, // sfix19_En18 
    input [18:0] Wgt_7_338, // sfix19_En18 
    input [18:0] Wgt_7_339, // sfix19_En18 
    input [18:0] Wgt_7_340, // sfix19_En18 
    input [18:0] Wgt_7_341, // sfix19_En18 
    input [18:0] Wgt_7_342, // sfix19_En18 
    input [18:0] Wgt_7_343, // sfix19_En18 
    input [18:0] Wgt_7_344, // sfix19_En18 
    input [18:0] Wgt_7_345, // sfix19_En18 
    input [18:0] Wgt_7_346, // sfix19_En18 
    input [18:0] Wgt_7_347, // sfix19_En18 
    input [18:0] Wgt_7_348, // sfix19_En18 
    input [18:0] Wgt_7_349, // sfix19_En18 
    input [18:0] Wgt_7_350, // sfix19_En18 
    input [18:0] Wgt_7_351, // sfix19_En18 
    input [18:0] Wgt_7_352, // sfix19_En18 
    input [18:0] Wgt_7_353, // sfix19_En18 
    input [18:0] Wgt_7_354, // sfix19_En18 
    input [18:0] Wgt_7_355, // sfix19_En18 
    input [18:0] Wgt_7_356, // sfix19_En18 
    input [18:0] Wgt_7_357, // sfix19_En18 
    input [18:0] Wgt_7_358, // sfix19_En18 
    input [18:0] Wgt_7_359, // sfix19_En18 
    input [18:0] Wgt_7_360, // sfix19_En18 
    input [18:0] Wgt_7_361, // sfix19_En18 
    input [18:0] Wgt_7_362, // sfix19_En18 
    input [18:0] Wgt_7_363, // sfix19_En18 
    input [18:0] Wgt_7_364, // sfix19_En18 
    input [18:0] Wgt_7_365, // sfix19_En18 
    input [18:0] Wgt_7_366, // sfix19_En18 
    input [18:0] Wgt_7_367, // sfix19_En18 
    input [18:0] Wgt_7_368, // sfix19_En18 
    input [18:0] Wgt_7_369, // sfix19_En18 
    input [18:0] Wgt_7_370, // sfix19_En18 
    input [18:0] Wgt_7_371, // sfix19_En18 
    input [18:0] Wgt_7_372, // sfix19_En18 
    input [18:0] Wgt_7_373, // sfix19_En18 
    input [18:0] Wgt_7_374, // sfix19_En18 
    input [18:0] Wgt_7_375, // sfix19_En18 
    input [18:0] Wgt_7_376, // sfix19_En18 
    input [18:0] Wgt_7_377, // sfix19_En18 
    input [18:0] Wgt_7_378, // sfix19_En18 
    input [18:0] Wgt_7_379, // sfix19_En18 
    input [18:0] Wgt_7_380, // sfix19_En18 
    input [18:0] Wgt_7_381, // sfix19_En18 
    input [18:0] Wgt_7_382, // sfix19_En18 
    input [18:0] Wgt_7_383, // sfix19_En18 
    input [18:0] Wgt_7_384, // sfix19_En18 
    input [18:0] Wgt_7_385, // sfix19_En18 
    input [18:0] Wgt_7_386, // sfix19_En18 
    input [18:0] Wgt_7_387, // sfix19_En18 
    input [18:0] Wgt_7_388, // sfix19_En18 
    input [18:0] Wgt_7_389, // sfix19_En18 
    input [18:0] Wgt_7_390, // sfix19_En18 
    input [18:0] Wgt_7_391, // sfix19_En18 
    input [18:0] Wgt_7_392, // sfix19_En18 
    input [18:0] Wgt_7_393, // sfix19_En18 
    input [18:0] Wgt_7_394, // sfix19_En18 
    input [18:0] Wgt_7_395, // sfix19_En18 
    input [18:0] Wgt_7_396, // sfix19_En18 
    input [18:0] Wgt_7_397, // sfix19_En18 
    input [18:0] Wgt_7_398, // sfix19_En18 
    input [18:0] Wgt_7_399, // sfix19_En18 
    input [18:0] Wgt_7_400, // sfix19_En18 
    input [18:0] Wgt_7_401, // sfix19_En18 
    input [18:0] Wgt_7_402, // sfix19_En18 
    input [18:0] Wgt_7_403, // sfix19_En18 
    input [18:0] Wgt_7_404, // sfix19_En18 
    input [18:0] Wgt_7_405, // sfix19_En18 
    input [18:0] Wgt_7_406, // sfix19_En18 
    input [18:0] Wgt_7_407, // sfix19_En18 
    input [18:0] Wgt_7_408, // sfix19_En18 
    input [18:0] Wgt_7_409, // sfix19_En18 
    input [18:0] Wgt_7_410, // sfix19_En18 
    input [18:0] Wgt_7_411, // sfix19_En18 
    input [18:0] Wgt_7_412, // sfix19_En18 
    input [18:0] Wgt_7_413, // sfix19_En18 
    input [18:0] Wgt_7_414, // sfix19_En18 
    input [18:0] Wgt_7_415, // sfix19_En18 
    input [18:0] Wgt_7_416, // sfix19_En18 
    input [18:0] Wgt_7_417, // sfix19_En18 
    input [18:0] Wgt_7_418, // sfix19_En18 
    input [18:0] Wgt_7_419, // sfix19_En18 
    input [18:0] Wgt_7_420, // sfix19_En18 
    input [18:0] Wgt_7_421, // sfix19_En18 
    input [18:0] Wgt_7_422, // sfix19_En18 
    input [18:0] Wgt_7_423, // sfix19_En18 
    input [18:0] Wgt_7_424, // sfix19_En18 
    input [18:0] Wgt_7_425, // sfix19_En18 
    input [18:0] Wgt_7_426, // sfix19_En18 
    input [18:0] Wgt_7_427, // sfix19_En18 
    input [18:0] Wgt_7_428, // sfix19_En18 
    input [18:0] Wgt_7_429, // sfix19_En18 
    input [18:0] Wgt_7_430, // sfix19_En18 
    input [18:0] Wgt_7_431, // sfix19_En18 
    input [18:0] Wgt_7_432, // sfix19_En18 
    input [18:0] Wgt_7_433, // sfix19_En18 
    input [18:0] Wgt_7_434, // sfix19_En18 
    input [18:0] Wgt_7_435, // sfix19_En18 
    input [18:0] Wgt_7_436, // sfix19_En18 
    input [18:0] Wgt_7_437, // sfix19_En18 
    input [18:0] Wgt_7_438, // sfix19_En18 
    input [18:0] Wgt_7_439, // sfix19_En18 
    input [18:0] Wgt_7_440, // sfix19_En18 
    input [18:0] Wgt_7_441, // sfix19_En18 
    input [18:0] Wgt_7_442, // sfix19_En18 
    input [18:0] Wgt_7_443, // sfix19_En18 
    input [18:0] Wgt_7_444, // sfix19_En18 
    input [18:0] Wgt_7_445, // sfix19_En18 
    input [18:0] Wgt_7_446, // sfix19_En18 
    input [18:0] Wgt_7_447, // sfix19_En18 
    input [18:0] Wgt_7_448, // sfix19_En18 
    input [18:0] Wgt_7_449, // sfix19_En18 
    input [18:0] Wgt_7_450, // sfix19_En18 
    input [18:0] Wgt_7_451, // sfix19_En18 
    input [18:0] Wgt_7_452, // sfix19_En18 
    input [18:0] Wgt_7_453, // sfix19_En18 
    input [18:0] Wgt_7_454, // sfix19_En18 
    input [18:0] Wgt_7_455, // sfix19_En18 
    input [18:0] Wgt_7_456, // sfix19_En18 
    input [18:0] Wgt_7_457, // sfix19_En18 
    input [18:0] Wgt_7_458, // sfix19_En18 
    input [18:0] Wgt_7_459, // sfix19_En18 
    input [18:0] Wgt_7_460, // sfix19_En18 
    input [18:0] Wgt_7_461, // sfix19_En18 
    input [18:0] Wgt_7_462, // sfix19_En18 
    input [18:0] Wgt_7_463, // sfix19_En18 
    input [18:0] Wgt_7_464, // sfix19_En18 
    input [18:0] Wgt_7_465, // sfix19_En18 
    input [18:0] Wgt_7_466, // sfix19_En18 
    input [18:0] Wgt_7_467, // sfix19_En18 
    input [18:0] Wgt_7_468, // sfix19_En18 
    input [18:0] Wgt_7_469, // sfix19_En18 
    input [18:0] Wgt_7_470, // sfix19_En18 
    input [18:0] Wgt_7_471, // sfix19_En18 
    input [18:0] Wgt_7_472, // sfix19_En18 
    input [18:0] Wgt_7_473, // sfix19_En18 
    input [18:0] Wgt_7_474, // sfix19_En18 
    input [18:0] Wgt_7_475, // sfix19_En18 
    input [18:0] Wgt_7_476, // sfix19_En18 
    input [18:0] Wgt_7_477, // sfix19_En18 
    input [18:0] Wgt_7_478, // sfix19_En18 
    input [18:0] Wgt_7_479, // sfix19_En18 
    input [18:0] Wgt_7_480, // sfix19_En18 
    input [18:0] Wgt_7_481, // sfix19_En18 
    input [18:0] Wgt_7_482, // sfix19_En18 
    input [18:0] Wgt_7_483, // sfix19_En18 
    input [18:0] Wgt_7_484, // sfix19_En18 
    input [18:0] Wgt_7_485, // sfix19_En18 
    input [18:0] Wgt_7_486, // sfix19_En18 
    input [18:0] Wgt_7_487, // sfix19_En18 
    input [18:0] Wgt_7_488, // sfix19_En18 
    input [18:0] Wgt_7_489, // sfix19_En18 
    input [18:0] Wgt_7_490, // sfix19_En18 
    input [18:0] Wgt_7_491, // sfix19_En18 
    input [18:0] Wgt_7_492, // sfix19_En18 
    input [18:0] Wgt_7_493, // sfix19_En18 
    input [18:0] Wgt_7_494, // sfix19_En18 
    input [18:0] Wgt_7_495, // sfix19_En18 
    input [18:0] Wgt_7_496, // sfix19_En18 
    input [18:0] Wgt_7_497, // sfix19_En18 
    input [18:0] Wgt_7_498, // sfix19_En18 
    input [18:0] Wgt_7_499, // sfix19_En18 
    input [18:0] Wgt_7_500, // sfix19_En18 
    input [18:0] Wgt_7_501, // sfix19_En18 
    input [18:0] Wgt_7_502, // sfix19_En18 
    input [18:0] Wgt_7_503, // sfix19_En18 
    input [18:0] Wgt_7_504, // sfix19_En18 
    input [18:0] Wgt_7_505, // sfix19_En18 
    input [18:0] Wgt_7_506, // sfix19_En18 
    input [18:0] Wgt_7_507, // sfix19_En18 
    input [18:0] Wgt_7_508, // sfix19_En18 
    input [18:0] Wgt_7_509, // sfix19_En18 
    input [18:0] Wgt_7_510, // sfix19_En18 
    input [18:0] Wgt_7_511, // sfix19_En18 
    input [18:0] Wgt_7_512, // sfix19_En18 
    input [18:0] Wgt_7_513, // sfix19_En18 
    input [18:0] Wgt_7_514, // sfix19_En18 
    input [18:0] Wgt_7_515, // sfix19_En18 
    input [18:0] Wgt_7_516, // sfix19_En18 
    input [18:0] Wgt_7_517, // sfix19_En18 
    input [18:0] Wgt_7_518, // sfix19_En18 
    input [18:0] Wgt_7_519, // sfix19_En18 
    input [18:0] Wgt_7_520, // sfix19_En18 
    input [18:0] Wgt_7_521, // sfix19_En18 
    input [18:0] Wgt_7_522, // sfix19_En18 
    input [18:0] Wgt_7_523, // sfix19_En18 
    input [18:0] Wgt_7_524, // sfix19_En18 
    input [18:0] Wgt_7_525, // sfix19_En18 
    input [18:0] Wgt_7_526, // sfix19_En18 
    input [18:0] Wgt_7_527, // sfix19_En18 
    input [18:0] Wgt_7_528, // sfix19_En18 
    input [18:0] Wgt_7_529, // sfix19_En18 
    input [18:0] Wgt_7_530, // sfix19_En18 
    input [18:0] Wgt_7_531, // sfix19_En18 
    input [18:0] Wgt_7_532, // sfix19_En18 
    input [18:0] Wgt_7_533, // sfix19_En18 
    input [18:0] Wgt_7_534, // sfix19_En18 
    input [18:0] Wgt_7_535, // sfix19_En18 
    input [18:0] Wgt_7_536, // sfix19_En18 
    input [18:0] Wgt_7_537, // sfix19_En18 
    input [18:0] Wgt_7_538, // sfix19_En18 
    input [18:0] Wgt_7_539, // sfix19_En18 
    input [18:0] Wgt_7_540, // sfix19_En18 
    input [18:0] Wgt_7_541, // sfix19_En18 
    input [18:0] Wgt_7_542, // sfix19_En18 
    input [18:0] Wgt_7_543, // sfix19_En18 
    input [18:0] Wgt_7_544, // sfix19_En18 
    input [18:0] Wgt_7_545, // sfix19_En18 
    input [18:0] Wgt_7_546, // sfix19_En18 
    input [18:0] Wgt_7_547, // sfix19_En18 
    input [18:0] Wgt_7_548, // sfix19_En18 
    input [18:0] Wgt_7_549, // sfix19_En18 
    input [18:0] Wgt_7_550, // sfix19_En18 
    input [18:0] Wgt_7_551, // sfix19_En18 
    input [18:0] Wgt_7_552, // sfix19_En18 
    input [18:0] Wgt_7_553, // sfix19_En18 
    input [18:0] Wgt_7_554, // sfix19_En18 
    input [18:0] Wgt_7_555, // sfix19_En18 
    input [18:0] Wgt_7_556, // sfix19_En18 
    input [18:0] Wgt_7_557, // sfix19_En18 
    input [18:0] Wgt_7_558, // sfix19_En18 
    input [18:0] Wgt_7_559, // sfix19_En18 
    input [18:0] Wgt_7_560, // sfix19_En18 
    input [18:0] Wgt_7_561, // sfix19_En18 
    input [18:0] Wgt_7_562, // sfix19_En18 
    input [18:0] Wgt_7_563, // sfix19_En18 
    input [18:0] Wgt_7_564, // sfix19_En18 
    input [18:0] Wgt_7_565, // sfix19_En18 
    input [18:0] Wgt_7_566, // sfix19_En18 
    input [18:0] Wgt_7_567, // sfix19_En18 
    input [18:0] Wgt_7_568, // sfix19_En18 
    input [18:0] Wgt_7_569, // sfix19_En18 
    input [18:0] Wgt_7_570, // sfix19_En18 
    input [18:0] Wgt_7_571, // sfix19_En18 
    input [18:0] Wgt_7_572, // sfix19_En18 
    input [18:0] Wgt_7_573, // sfix19_En18 
    input [18:0] Wgt_7_574, // sfix19_En18 
    input [18:0] Wgt_7_575, // sfix19_En18 
    input [18:0] Wgt_7_576, // sfix19_En18 
    input [18:0] Wgt_7_577, // sfix19_En18 
    input [18:0] Wgt_7_578, // sfix19_En18 
    input [18:0] Wgt_7_579, // sfix19_En18 
    input [18:0] Wgt_7_580, // sfix19_En18 
    input [18:0] Wgt_7_581, // sfix19_En18 
    input [18:0] Wgt_7_582, // sfix19_En18 
    input [18:0] Wgt_7_583, // sfix19_En18 
    input [18:0] Wgt_7_584, // sfix19_En18 
    input [18:0] Wgt_7_585, // sfix19_En18 
    input [18:0] Wgt_7_586, // sfix19_En18 
    input [18:0] Wgt_7_587, // sfix19_En18 
    input [18:0] Wgt_7_588, // sfix19_En18 
    input [18:0] Wgt_7_589, // sfix19_En18 
    input [18:0] Wgt_7_590, // sfix19_En18 
    input [18:0] Wgt_7_591, // sfix19_En18 
    input [18:0] Wgt_7_592, // sfix19_En18 
    input [18:0] Wgt_7_593, // sfix19_En18 
    input [18:0] Wgt_7_594, // sfix19_En18 
    input [18:0] Wgt_7_595, // sfix19_En18 
    input [18:0] Wgt_7_596, // sfix19_En18 
    input [18:0] Wgt_7_597, // sfix19_En18 
    input [18:0] Wgt_7_598, // sfix19_En18 
    input [18:0] Wgt_7_599, // sfix19_En18 
    input [18:0] Wgt_7_600, // sfix19_En18 
    input [18:0] Wgt_7_601, // sfix19_En18 
    input [18:0] Wgt_7_602, // sfix19_En18 
    input [18:0] Wgt_7_603, // sfix19_En18 
    input [18:0] Wgt_7_604, // sfix19_En18 
    input [18:0] Wgt_7_605, // sfix19_En18 
    input [18:0] Wgt_7_606, // sfix19_En18 
    input [18:0] Wgt_7_607, // sfix19_En18 
    input [18:0] Wgt_7_608, // sfix19_En18 
    input [18:0] Wgt_7_609, // sfix19_En18 
    input [18:0] Wgt_7_610, // sfix19_En18 
    input [18:0] Wgt_7_611, // sfix19_En18 
    input [18:0] Wgt_7_612, // sfix19_En18 
    input [18:0] Wgt_7_613, // sfix19_En18 
    input [18:0] Wgt_7_614, // sfix19_En18 
    input [18:0] Wgt_7_615, // sfix19_En18 
    input [18:0] Wgt_7_616, // sfix19_En18 
    input [18:0] Wgt_7_617, // sfix19_En18 
    input [18:0] Wgt_7_618, // sfix19_En18 
    input [18:0] Wgt_7_619, // sfix19_En18 
    input [18:0] Wgt_7_620, // sfix19_En18 
    input [18:0] Wgt_7_621, // sfix19_En18 
    input [18:0] Wgt_7_622, // sfix19_En18 
    input [18:0] Wgt_7_623, // sfix19_En18 
    input [18:0] Wgt_7_624, // sfix19_En18 
    input [18:0] Wgt_7_625, // sfix19_En18 
    input [18:0] Wgt_7_626, // sfix19_En18 
    input [18:0] Wgt_7_627, // sfix19_En18 
    input [18:0] Wgt_7_628, // sfix19_En18 
    input [18:0] Wgt_7_629, // sfix19_En18 
    input [18:0] Wgt_7_630, // sfix19_En18 
    input [18:0] Wgt_7_631, // sfix19_En18 
    input [18:0] Wgt_7_632, // sfix19_En18 
    input [18:0] Wgt_7_633, // sfix19_En18 
    input [18:0] Wgt_7_634, // sfix19_En18 
    input [18:0] Wgt_7_635, // sfix19_En18 
    input [18:0] Wgt_7_636, // sfix19_En18 
    input [18:0] Wgt_7_637, // sfix19_En18 
    input [18:0] Wgt_7_638, // sfix19_En18 
    input [18:0] Wgt_7_639, // sfix19_En18 
    input [18:0] Wgt_7_640, // sfix19_En18 
    input [18:0] Wgt_7_641, // sfix19_En18 
    input [18:0] Wgt_7_642, // sfix19_En18 
    input [18:0] Wgt_7_643, // sfix19_En18 
    input [18:0] Wgt_7_644, // sfix19_En18 
    input [18:0] Wgt_7_645, // sfix19_En18 
    input [18:0] Wgt_7_646, // sfix19_En18 
    input [18:0] Wgt_7_647, // sfix19_En18 
    input [18:0] Wgt_7_648, // sfix19_En18 
    input [18:0] Wgt_7_649, // sfix19_En18 
    input [18:0] Wgt_7_650, // sfix19_En18 
    input [18:0] Wgt_7_651, // sfix19_En18 
    input [18:0] Wgt_7_652, // sfix19_En18 
    input [18:0] Wgt_7_653, // sfix19_En18 
    input [18:0] Wgt_7_654, // sfix19_En18 
    input [18:0] Wgt_7_655, // sfix19_En18 
    input [18:0] Wgt_7_656, // sfix19_En18 
    input [18:0] Wgt_7_657, // sfix19_En18 
    input [18:0] Wgt_7_658, // sfix19_En18 
    input [18:0] Wgt_7_659, // sfix19_En18 
    input [18:0] Wgt_7_660, // sfix19_En18 
    input [18:0] Wgt_7_661, // sfix19_En18 
    input [18:0] Wgt_7_662, // sfix19_En18 
    input [18:0] Wgt_7_663, // sfix19_En18 
    input [18:0] Wgt_7_664, // sfix19_En18 
    input [18:0] Wgt_7_665, // sfix19_En18 
    input [18:0] Wgt_7_666, // sfix19_En18 
    input [18:0] Wgt_7_667, // sfix19_En18 
    input [18:0] Wgt_7_668, // sfix19_En18 
    input [18:0] Wgt_7_669, // sfix19_En18 
    input [18:0] Wgt_7_670, // sfix19_En18 
    input [18:0] Wgt_7_671, // sfix19_En18 
    input [18:0] Wgt_7_672, // sfix19_En18 
    input [18:0] Wgt_7_673, // sfix19_En18 
    input [18:0] Wgt_7_674, // sfix19_En18 
    input [18:0] Wgt_7_675, // sfix19_En18 
    input [18:0] Wgt_7_676, // sfix19_En18 
    input [18:0] Wgt_7_677, // sfix19_En18 
    input [18:0] Wgt_7_678, // sfix19_En18 
    input [18:0] Wgt_7_679, // sfix19_En18 
    input [18:0] Wgt_7_680, // sfix19_En18 
    input [18:0] Wgt_7_681, // sfix19_En18 
    input [18:0] Wgt_7_682, // sfix19_En18 
    input [18:0] Wgt_7_683, // sfix19_En18 
    input [18:0] Wgt_7_684, // sfix19_En18 
    input [18:0] Wgt_7_685, // sfix19_En18 
    input [18:0] Wgt_7_686, // sfix19_En18 
    input [18:0] Wgt_7_687, // sfix19_En18 
    input [18:0] Wgt_7_688, // sfix19_En18 
    input [18:0] Wgt_7_689, // sfix19_En18 
    input [18:0] Wgt_7_690, // sfix19_En18 
    input [18:0] Wgt_7_691, // sfix19_En18 
    input [18:0] Wgt_7_692, // sfix19_En18 
    input [18:0] Wgt_7_693, // sfix19_En18 
    input [18:0] Wgt_7_694, // sfix19_En18 
    input [18:0] Wgt_7_695, // sfix19_En18 
    input [18:0] Wgt_7_696, // sfix19_En18 
    input [18:0] Wgt_7_697, // sfix19_En18 
    input [18:0] Wgt_7_698, // sfix19_En18 
    input [18:0] Wgt_7_699, // sfix19_En18 
    input [18:0] Wgt_7_700, // sfix19_En18 
    input [18:0] Wgt_7_701, // sfix19_En18 
    input [18:0] Wgt_7_702, // sfix19_En18 
    input [18:0] Wgt_7_703, // sfix19_En18 
    input [18:0] Wgt_7_704, // sfix19_En18 
    input [18:0] Wgt_7_705, // sfix19_En18 
    input [18:0] Wgt_7_706, // sfix19_En18 
    input [18:0] Wgt_7_707, // sfix19_En18 
    input [18:0] Wgt_7_708, // sfix19_En18 
    input [18:0] Wgt_7_709, // sfix19_En18 
    input [18:0] Wgt_7_710, // sfix19_En18 
    input [18:0] Wgt_7_711, // sfix19_En18 
    input [18:0] Wgt_7_712, // sfix19_En18 
    input [18:0] Wgt_7_713, // sfix19_En18 
    input [18:0] Wgt_7_714, // sfix19_En18 
    input [18:0] Wgt_7_715, // sfix19_En18 
    input [18:0] Wgt_7_716, // sfix19_En18 
    input [18:0] Wgt_7_717, // sfix19_En18 
    input [18:0] Wgt_7_718, // sfix19_En18 
    input [18:0] Wgt_7_719, // sfix19_En18 
    input [18:0] Wgt_7_720, // sfix19_En18 
    input [18:0] Wgt_7_721, // sfix19_En18 
    input [18:0] Wgt_7_722, // sfix19_En18 
    input [18:0] Wgt_7_723, // sfix19_En18 
    input [18:0] Wgt_7_724, // sfix19_En18 
    input [18:0] Wgt_7_725, // sfix19_En18 
    input [18:0] Wgt_7_726, // sfix19_En18 
    input [18:0] Wgt_7_727, // sfix19_En18 
    input [18:0] Wgt_7_728, // sfix19_En18 
    input [18:0] Wgt_7_729, // sfix19_En18 
    input [18:0] Wgt_7_730, // sfix19_En18 
    input [18:0] Wgt_7_731, // sfix19_En18 
    input [18:0] Wgt_7_732, // sfix19_En18 
    input [18:0] Wgt_7_733, // sfix19_En18 
    input [18:0] Wgt_7_734, // sfix19_En18 
    input [18:0] Wgt_7_735, // sfix19_En18 
    input [18:0] Wgt_7_736, // sfix19_En18 
    input [18:0] Wgt_7_737, // sfix19_En18 
    input [18:0] Wgt_7_738, // sfix19_En18 
    input [18:0] Wgt_7_739, // sfix19_En18 
    input [18:0] Wgt_7_740, // sfix19_En18 
    input [18:0] Wgt_7_741, // sfix19_En18 
    input [18:0] Wgt_7_742, // sfix19_En18 
    input [18:0] Wgt_7_743, // sfix19_En18 
    input [18:0] Wgt_7_744, // sfix19_En18 
    input [18:0] Wgt_7_745, // sfix19_En18 
    input [18:0] Wgt_7_746, // sfix19_En18 
    input [18:0] Wgt_7_747, // sfix19_En18 
    input [18:0] Wgt_7_748, // sfix19_En18 
    input [18:0] Wgt_7_749, // sfix19_En18 
    input [18:0] Wgt_7_750, // sfix19_En18 
    input [18:0] Wgt_7_751, // sfix19_En18 
    input [18:0] Wgt_7_752, // sfix19_En18 
    input [18:0] Wgt_7_753, // sfix19_En18 
    input [18:0] Wgt_7_754, // sfix19_En18 
    input [18:0] Wgt_7_755, // sfix19_En18 
    input [18:0] Wgt_7_756, // sfix19_En18 
    input [18:0] Wgt_7_757, // sfix19_En18 
    input [18:0] Wgt_7_758, // sfix19_En18 
    input [18:0] Wgt_7_759, // sfix19_En18 
    input [18:0] Wgt_7_760, // sfix19_En18 
    input [18:0] Wgt_7_761, // sfix19_En18 
    input [18:0] Wgt_7_762, // sfix19_En18 
    input [18:0] Wgt_7_763, // sfix19_En18 
    input [18:0] Wgt_7_764, // sfix19_En18 
    input [18:0] Wgt_7_765, // sfix19_En18 
    input [18:0] Wgt_7_766, // sfix19_En18 
    input [18:0] Wgt_7_767, // sfix19_En18 
    input [18:0] Wgt_7_768, // sfix19_En18 
    input [18:0] Wgt_7_769, // sfix19_En18 
    input [18:0] Wgt_7_770, // sfix19_En18 
    input [18:0] Wgt_7_771, // sfix19_En18 
    input [18:0] Wgt_7_772, // sfix19_En18 
    input [18:0] Wgt_7_773, // sfix19_En18 
    input [18:0] Wgt_7_774, // sfix19_En18 
    input [18:0] Wgt_7_775, // sfix19_En18 
    input [18:0] Wgt_7_776, // sfix19_En18 
    input [18:0] Wgt_7_777, // sfix19_En18 
    input [18:0] Wgt_7_778, // sfix19_En18 
    input [18:0] Wgt_7_779, // sfix19_En18 
    input [18:0] Wgt_7_780, // sfix19_En18 
    input [18:0] Wgt_7_781, // sfix19_En18 
    input [18:0] Wgt_7_782, // sfix19_En18 
    input [18:0] Wgt_7_783, // sfix19_En18 
    input [18:0] Wgt_7_784, // sfix19_En18 
    input [18:0] Wgt_8_0, // sfix19_En18 
    input [18:0] Wgt_8_1, // sfix19_En18 
    input [18:0] Wgt_8_2, // sfix19_En18 
    input [18:0] Wgt_8_3, // sfix19_En18 
    input [18:0] Wgt_8_4, // sfix19_En18 
    input [18:0] Wgt_8_5, // sfix19_En18 
    input [18:0] Wgt_8_6, // sfix19_En18 
    input [18:0] Wgt_8_7, // sfix19_En18 
    input [18:0] Wgt_8_8, // sfix19_En18 
    input [18:0] Wgt_8_9, // sfix19_En18 
    input [18:0] Wgt_8_10, // sfix19_En18 
    input [18:0] Wgt_8_11, // sfix19_En18 
    input [18:0] Wgt_8_12, // sfix19_En18 
    input [18:0] Wgt_8_13, // sfix19_En18 
    input [18:0] Wgt_8_14, // sfix19_En18 
    input [18:0] Wgt_8_15, // sfix19_En18 
    input [18:0] Wgt_8_16, // sfix19_En18 
    input [18:0] Wgt_8_17, // sfix19_En18 
    input [18:0] Wgt_8_18, // sfix19_En18 
    input [18:0] Wgt_8_19, // sfix19_En18 
    input [18:0] Wgt_8_20, // sfix19_En18 
    input [18:0] Wgt_8_21, // sfix19_En18 
    input [18:0] Wgt_8_22, // sfix19_En18 
    input [18:0] Wgt_8_23, // sfix19_En18 
    input [18:0] Wgt_8_24, // sfix19_En18 
    input [18:0] Wgt_8_25, // sfix19_En18 
    input [18:0] Wgt_8_26, // sfix19_En18 
    input [18:0] Wgt_8_27, // sfix19_En18 
    input [18:0] Wgt_8_28, // sfix19_En18 
    input [18:0] Wgt_8_29, // sfix19_En18 
    input [18:0] Wgt_8_30, // sfix19_En18 
    input [18:0] Wgt_8_31, // sfix19_En18 
    input [18:0] Wgt_8_32, // sfix19_En18 
    input [18:0] Wgt_8_33, // sfix19_En18 
    input [18:0] Wgt_8_34, // sfix19_En18 
    input [18:0] Wgt_8_35, // sfix19_En18 
    input [18:0] Wgt_8_36, // sfix19_En18 
    input [18:0] Wgt_8_37, // sfix19_En18 
    input [18:0] Wgt_8_38, // sfix19_En18 
    input [18:0] Wgt_8_39, // sfix19_En18 
    input [18:0] Wgt_8_40, // sfix19_En18 
    input [18:0] Wgt_8_41, // sfix19_En18 
    input [18:0] Wgt_8_42, // sfix19_En18 
    input [18:0] Wgt_8_43, // sfix19_En18 
    input [18:0] Wgt_8_44, // sfix19_En18 
    input [18:0] Wgt_8_45, // sfix19_En18 
    input [18:0] Wgt_8_46, // sfix19_En18 
    input [18:0] Wgt_8_47, // sfix19_En18 
    input [18:0] Wgt_8_48, // sfix19_En18 
    input [18:0] Wgt_8_49, // sfix19_En18 
    input [18:0] Wgt_8_50, // sfix19_En18 
    input [18:0] Wgt_8_51, // sfix19_En18 
    input [18:0] Wgt_8_52, // sfix19_En18 
    input [18:0] Wgt_8_53, // sfix19_En18 
    input [18:0] Wgt_8_54, // sfix19_En18 
    input [18:0] Wgt_8_55, // sfix19_En18 
    input [18:0] Wgt_8_56, // sfix19_En18 
    input [18:0] Wgt_8_57, // sfix19_En18 
    input [18:0] Wgt_8_58, // sfix19_En18 
    input [18:0] Wgt_8_59, // sfix19_En18 
    input [18:0] Wgt_8_60, // sfix19_En18 
    input [18:0] Wgt_8_61, // sfix19_En18 
    input [18:0] Wgt_8_62, // sfix19_En18 
    input [18:0] Wgt_8_63, // sfix19_En18 
    input [18:0] Wgt_8_64, // sfix19_En18 
    input [18:0] Wgt_8_65, // sfix19_En18 
    input [18:0] Wgt_8_66, // sfix19_En18 
    input [18:0] Wgt_8_67, // sfix19_En18 
    input [18:0] Wgt_8_68, // sfix19_En18 
    input [18:0] Wgt_8_69, // sfix19_En18 
    input [18:0] Wgt_8_70, // sfix19_En18 
    input [18:0] Wgt_8_71, // sfix19_En18 
    input [18:0] Wgt_8_72, // sfix19_En18 
    input [18:0] Wgt_8_73, // sfix19_En18 
    input [18:0] Wgt_8_74, // sfix19_En18 
    input [18:0] Wgt_8_75, // sfix19_En18 
    input [18:0] Wgt_8_76, // sfix19_En18 
    input [18:0] Wgt_8_77, // sfix19_En18 
    input [18:0] Wgt_8_78, // sfix19_En18 
    input [18:0] Wgt_8_79, // sfix19_En18 
    input [18:0] Wgt_8_80, // sfix19_En18 
    input [18:0] Wgt_8_81, // sfix19_En18 
    input [18:0] Wgt_8_82, // sfix19_En18 
    input [18:0] Wgt_8_83, // sfix19_En18 
    input [18:0] Wgt_8_84, // sfix19_En18 
    input [18:0] Wgt_8_85, // sfix19_En18 
    input [18:0] Wgt_8_86, // sfix19_En18 
    input [18:0] Wgt_8_87, // sfix19_En18 
    input [18:0] Wgt_8_88, // sfix19_En18 
    input [18:0] Wgt_8_89, // sfix19_En18 
    input [18:0] Wgt_8_90, // sfix19_En18 
    input [18:0] Wgt_8_91, // sfix19_En18 
    input [18:0] Wgt_8_92, // sfix19_En18 
    input [18:0] Wgt_8_93, // sfix19_En18 
    input [18:0] Wgt_8_94, // sfix19_En18 
    input [18:0] Wgt_8_95, // sfix19_En18 
    input [18:0] Wgt_8_96, // sfix19_En18 
    input [18:0] Wgt_8_97, // sfix19_En18 
    input [18:0] Wgt_8_98, // sfix19_En18 
    input [18:0] Wgt_8_99, // sfix19_En18 
    input [18:0] Wgt_8_100, // sfix19_En18 
    input [18:0] Wgt_8_101, // sfix19_En18 
    input [18:0] Wgt_8_102, // sfix19_En18 
    input [18:0] Wgt_8_103, // sfix19_En18 
    input [18:0] Wgt_8_104, // sfix19_En18 
    input [18:0] Wgt_8_105, // sfix19_En18 
    input [18:0] Wgt_8_106, // sfix19_En18 
    input [18:0] Wgt_8_107, // sfix19_En18 
    input [18:0] Wgt_8_108, // sfix19_En18 
    input [18:0] Wgt_8_109, // sfix19_En18 
    input [18:0] Wgt_8_110, // sfix19_En18 
    input [18:0] Wgt_8_111, // sfix19_En18 
    input [18:0] Wgt_8_112, // sfix19_En18 
    input [18:0] Wgt_8_113, // sfix19_En18 
    input [18:0] Wgt_8_114, // sfix19_En18 
    input [18:0] Wgt_8_115, // sfix19_En18 
    input [18:0] Wgt_8_116, // sfix19_En18 
    input [18:0] Wgt_8_117, // sfix19_En18 
    input [18:0] Wgt_8_118, // sfix19_En18 
    input [18:0] Wgt_8_119, // sfix19_En18 
    input [18:0] Wgt_8_120, // sfix19_En18 
    input [18:0] Wgt_8_121, // sfix19_En18 
    input [18:0] Wgt_8_122, // sfix19_En18 
    input [18:0] Wgt_8_123, // sfix19_En18 
    input [18:0] Wgt_8_124, // sfix19_En18 
    input [18:0] Wgt_8_125, // sfix19_En18 
    input [18:0] Wgt_8_126, // sfix19_En18 
    input [18:0] Wgt_8_127, // sfix19_En18 
    input [18:0] Wgt_8_128, // sfix19_En18 
    input [18:0] Wgt_8_129, // sfix19_En18 
    input [18:0] Wgt_8_130, // sfix19_En18 
    input [18:0] Wgt_8_131, // sfix19_En18 
    input [18:0] Wgt_8_132, // sfix19_En18 
    input [18:0] Wgt_8_133, // sfix19_En18 
    input [18:0] Wgt_8_134, // sfix19_En18 
    input [18:0] Wgt_8_135, // sfix19_En18 
    input [18:0] Wgt_8_136, // sfix19_En18 
    input [18:0] Wgt_8_137, // sfix19_En18 
    input [18:0] Wgt_8_138, // sfix19_En18 
    input [18:0] Wgt_8_139, // sfix19_En18 
    input [18:0] Wgt_8_140, // sfix19_En18 
    input [18:0] Wgt_8_141, // sfix19_En18 
    input [18:0] Wgt_8_142, // sfix19_En18 
    input [18:0] Wgt_8_143, // sfix19_En18 
    input [18:0] Wgt_8_144, // sfix19_En18 
    input [18:0] Wgt_8_145, // sfix19_En18 
    input [18:0] Wgt_8_146, // sfix19_En18 
    input [18:0] Wgt_8_147, // sfix19_En18 
    input [18:0] Wgt_8_148, // sfix19_En18 
    input [18:0] Wgt_8_149, // sfix19_En18 
    input [18:0] Wgt_8_150, // sfix19_En18 
    input [18:0] Wgt_8_151, // sfix19_En18 
    input [18:0] Wgt_8_152, // sfix19_En18 
    input [18:0] Wgt_8_153, // sfix19_En18 
    input [18:0] Wgt_8_154, // sfix19_En18 
    input [18:0] Wgt_8_155, // sfix19_En18 
    input [18:0] Wgt_8_156, // sfix19_En18 
    input [18:0] Wgt_8_157, // sfix19_En18 
    input [18:0] Wgt_8_158, // sfix19_En18 
    input [18:0] Wgt_8_159, // sfix19_En18 
    input [18:0] Wgt_8_160, // sfix19_En18 
    input [18:0] Wgt_8_161, // sfix19_En18 
    input [18:0] Wgt_8_162, // sfix19_En18 
    input [18:0] Wgt_8_163, // sfix19_En18 
    input [18:0] Wgt_8_164, // sfix19_En18 
    input [18:0] Wgt_8_165, // sfix19_En18 
    input [18:0] Wgt_8_166, // sfix19_En18 
    input [18:0] Wgt_8_167, // sfix19_En18 
    input [18:0] Wgt_8_168, // sfix19_En18 
    input [18:0] Wgt_8_169, // sfix19_En18 
    input [18:0] Wgt_8_170, // sfix19_En18 
    input [18:0] Wgt_8_171, // sfix19_En18 
    input [18:0] Wgt_8_172, // sfix19_En18 
    input [18:0] Wgt_8_173, // sfix19_En18 
    input [18:0] Wgt_8_174, // sfix19_En18 
    input [18:0] Wgt_8_175, // sfix19_En18 
    input [18:0] Wgt_8_176, // sfix19_En18 
    input [18:0] Wgt_8_177, // sfix19_En18 
    input [18:0] Wgt_8_178, // sfix19_En18 
    input [18:0] Wgt_8_179, // sfix19_En18 
    input [18:0] Wgt_8_180, // sfix19_En18 
    input [18:0] Wgt_8_181, // sfix19_En18 
    input [18:0] Wgt_8_182, // sfix19_En18 
    input [18:0] Wgt_8_183, // sfix19_En18 
    input [18:0] Wgt_8_184, // sfix19_En18 
    input [18:0] Wgt_8_185, // sfix19_En18 
    input [18:0] Wgt_8_186, // sfix19_En18 
    input [18:0] Wgt_8_187, // sfix19_En18 
    input [18:0] Wgt_8_188, // sfix19_En18 
    input [18:0] Wgt_8_189, // sfix19_En18 
    input [18:0] Wgt_8_190, // sfix19_En18 
    input [18:0] Wgt_8_191, // sfix19_En18 
    input [18:0] Wgt_8_192, // sfix19_En18 
    input [18:0] Wgt_8_193, // sfix19_En18 
    input [18:0] Wgt_8_194, // sfix19_En18 
    input [18:0] Wgt_8_195, // sfix19_En18 
    input [18:0] Wgt_8_196, // sfix19_En18 
    input [18:0] Wgt_8_197, // sfix19_En18 
    input [18:0] Wgt_8_198, // sfix19_En18 
    input [18:0] Wgt_8_199, // sfix19_En18 
    input [18:0] Wgt_8_200, // sfix19_En18 
    input [18:0] Wgt_8_201, // sfix19_En18 
    input [18:0] Wgt_8_202, // sfix19_En18 
    input [18:0] Wgt_8_203, // sfix19_En18 
    input [18:0] Wgt_8_204, // sfix19_En18 
    input [18:0] Wgt_8_205, // sfix19_En18 
    input [18:0] Wgt_8_206, // sfix19_En18 
    input [18:0] Wgt_8_207, // sfix19_En18 
    input [18:0] Wgt_8_208, // sfix19_En18 
    input [18:0] Wgt_8_209, // sfix19_En18 
    input [18:0] Wgt_8_210, // sfix19_En18 
    input [18:0] Wgt_8_211, // sfix19_En18 
    input [18:0] Wgt_8_212, // sfix19_En18 
    input [18:0] Wgt_8_213, // sfix19_En18 
    input [18:0] Wgt_8_214, // sfix19_En18 
    input [18:0] Wgt_8_215, // sfix19_En18 
    input [18:0] Wgt_8_216, // sfix19_En18 
    input [18:0] Wgt_8_217, // sfix19_En18 
    input [18:0] Wgt_8_218, // sfix19_En18 
    input [18:0] Wgt_8_219, // sfix19_En18 
    input [18:0] Wgt_8_220, // sfix19_En18 
    input [18:0] Wgt_8_221, // sfix19_En18 
    input [18:0] Wgt_8_222, // sfix19_En18 
    input [18:0] Wgt_8_223, // sfix19_En18 
    input [18:0] Wgt_8_224, // sfix19_En18 
    input [18:0] Wgt_8_225, // sfix19_En18 
    input [18:0] Wgt_8_226, // sfix19_En18 
    input [18:0] Wgt_8_227, // sfix19_En18 
    input [18:0] Wgt_8_228, // sfix19_En18 
    input [18:0] Wgt_8_229, // sfix19_En18 
    input [18:0] Wgt_8_230, // sfix19_En18 
    input [18:0] Wgt_8_231, // sfix19_En18 
    input [18:0] Wgt_8_232, // sfix19_En18 
    input [18:0] Wgt_8_233, // sfix19_En18 
    input [18:0] Wgt_8_234, // sfix19_En18 
    input [18:0] Wgt_8_235, // sfix19_En18 
    input [18:0] Wgt_8_236, // sfix19_En18 
    input [18:0] Wgt_8_237, // sfix19_En18 
    input [18:0] Wgt_8_238, // sfix19_En18 
    input [18:0] Wgt_8_239, // sfix19_En18 
    input [18:0] Wgt_8_240, // sfix19_En18 
    input [18:0] Wgt_8_241, // sfix19_En18 
    input [18:0] Wgt_8_242, // sfix19_En18 
    input [18:0] Wgt_8_243, // sfix19_En18 
    input [18:0] Wgt_8_244, // sfix19_En18 
    input [18:0] Wgt_8_245, // sfix19_En18 
    input [18:0] Wgt_8_246, // sfix19_En18 
    input [18:0] Wgt_8_247, // sfix19_En18 
    input [18:0] Wgt_8_248, // sfix19_En18 
    input [18:0] Wgt_8_249, // sfix19_En18 
    input [18:0] Wgt_8_250, // sfix19_En18 
    input [18:0] Wgt_8_251, // sfix19_En18 
    input [18:0] Wgt_8_252, // sfix19_En18 
    input [18:0] Wgt_8_253, // sfix19_En18 
    input [18:0] Wgt_8_254, // sfix19_En18 
    input [18:0] Wgt_8_255, // sfix19_En18 
    input [18:0] Wgt_8_256, // sfix19_En18 
    input [18:0] Wgt_8_257, // sfix19_En18 
    input [18:0] Wgt_8_258, // sfix19_En18 
    input [18:0] Wgt_8_259, // sfix19_En18 
    input [18:0] Wgt_8_260, // sfix19_En18 
    input [18:0] Wgt_8_261, // sfix19_En18 
    input [18:0] Wgt_8_262, // sfix19_En18 
    input [18:0] Wgt_8_263, // sfix19_En18 
    input [18:0] Wgt_8_264, // sfix19_En18 
    input [18:0] Wgt_8_265, // sfix19_En18 
    input [18:0] Wgt_8_266, // sfix19_En18 
    input [18:0] Wgt_8_267, // sfix19_En18 
    input [18:0] Wgt_8_268, // sfix19_En18 
    input [18:0] Wgt_8_269, // sfix19_En18 
    input [18:0] Wgt_8_270, // sfix19_En18 
    input [18:0] Wgt_8_271, // sfix19_En18 
    input [18:0] Wgt_8_272, // sfix19_En18 
    input [18:0] Wgt_8_273, // sfix19_En18 
    input [18:0] Wgt_8_274, // sfix19_En18 
    input [18:0] Wgt_8_275, // sfix19_En18 
    input [18:0] Wgt_8_276, // sfix19_En18 
    input [18:0] Wgt_8_277, // sfix19_En18 
    input [18:0] Wgt_8_278, // sfix19_En18 
    input [18:0] Wgt_8_279, // sfix19_En18 
    input [18:0] Wgt_8_280, // sfix19_En18 
    input [18:0] Wgt_8_281, // sfix19_En18 
    input [18:0] Wgt_8_282, // sfix19_En18 
    input [18:0] Wgt_8_283, // sfix19_En18 
    input [18:0] Wgt_8_284, // sfix19_En18 
    input [18:0] Wgt_8_285, // sfix19_En18 
    input [18:0] Wgt_8_286, // sfix19_En18 
    input [18:0] Wgt_8_287, // sfix19_En18 
    input [18:0] Wgt_8_288, // sfix19_En18 
    input [18:0] Wgt_8_289, // sfix19_En18 
    input [18:0] Wgt_8_290, // sfix19_En18 
    input [18:0] Wgt_8_291, // sfix19_En18 
    input [18:0] Wgt_8_292, // sfix19_En18 
    input [18:0] Wgt_8_293, // sfix19_En18 
    input [18:0] Wgt_8_294, // sfix19_En18 
    input [18:0] Wgt_8_295, // sfix19_En18 
    input [18:0] Wgt_8_296, // sfix19_En18 
    input [18:0] Wgt_8_297, // sfix19_En18 
    input [18:0] Wgt_8_298, // sfix19_En18 
    input [18:0] Wgt_8_299, // sfix19_En18 
    input [18:0] Wgt_8_300, // sfix19_En18 
    input [18:0] Wgt_8_301, // sfix19_En18 
    input [18:0] Wgt_8_302, // sfix19_En18 
    input [18:0] Wgt_8_303, // sfix19_En18 
    input [18:0] Wgt_8_304, // sfix19_En18 
    input [18:0] Wgt_8_305, // sfix19_En18 
    input [18:0] Wgt_8_306, // sfix19_En18 
    input [18:0] Wgt_8_307, // sfix19_En18 
    input [18:0] Wgt_8_308, // sfix19_En18 
    input [18:0] Wgt_8_309, // sfix19_En18 
    input [18:0] Wgt_8_310, // sfix19_En18 
    input [18:0] Wgt_8_311, // sfix19_En18 
    input [18:0] Wgt_8_312, // sfix19_En18 
    input [18:0] Wgt_8_313, // sfix19_En18 
    input [18:0] Wgt_8_314, // sfix19_En18 
    input [18:0] Wgt_8_315, // sfix19_En18 
    input [18:0] Wgt_8_316, // sfix19_En18 
    input [18:0] Wgt_8_317, // sfix19_En18 
    input [18:0] Wgt_8_318, // sfix19_En18 
    input [18:0] Wgt_8_319, // sfix19_En18 
    input [18:0] Wgt_8_320, // sfix19_En18 
    input [18:0] Wgt_8_321, // sfix19_En18 
    input [18:0] Wgt_8_322, // sfix19_En18 
    input [18:0] Wgt_8_323, // sfix19_En18 
    input [18:0] Wgt_8_324, // sfix19_En18 
    input [18:0] Wgt_8_325, // sfix19_En18 
    input [18:0] Wgt_8_326, // sfix19_En18 
    input [18:0] Wgt_8_327, // sfix19_En18 
    input [18:0] Wgt_8_328, // sfix19_En18 
    input [18:0] Wgt_8_329, // sfix19_En18 
    input [18:0] Wgt_8_330, // sfix19_En18 
    input [18:0] Wgt_8_331, // sfix19_En18 
    input [18:0] Wgt_8_332, // sfix19_En18 
    input [18:0] Wgt_8_333, // sfix19_En18 
    input [18:0] Wgt_8_334, // sfix19_En18 
    input [18:0] Wgt_8_335, // sfix19_En18 
    input [18:0] Wgt_8_336, // sfix19_En18 
    input [18:0] Wgt_8_337, // sfix19_En18 
    input [18:0] Wgt_8_338, // sfix19_En18 
    input [18:0] Wgt_8_339, // sfix19_En18 
    input [18:0] Wgt_8_340, // sfix19_En18 
    input [18:0] Wgt_8_341, // sfix19_En18 
    input [18:0] Wgt_8_342, // sfix19_En18 
    input [18:0] Wgt_8_343, // sfix19_En18 
    input [18:0] Wgt_8_344, // sfix19_En18 
    input [18:0] Wgt_8_345, // sfix19_En18 
    input [18:0] Wgt_8_346, // sfix19_En18 
    input [18:0] Wgt_8_347, // sfix19_En18 
    input [18:0] Wgt_8_348, // sfix19_En18 
    input [18:0] Wgt_8_349, // sfix19_En18 
    input [18:0] Wgt_8_350, // sfix19_En18 
    input [18:0] Wgt_8_351, // sfix19_En18 
    input [18:0] Wgt_8_352, // sfix19_En18 
    input [18:0] Wgt_8_353, // sfix19_En18 
    input [18:0] Wgt_8_354, // sfix19_En18 
    input [18:0] Wgt_8_355, // sfix19_En18 
    input [18:0] Wgt_8_356, // sfix19_En18 
    input [18:0] Wgt_8_357, // sfix19_En18 
    input [18:0] Wgt_8_358, // sfix19_En18 
    input [18:0] Wgt_8_359, // sfix19_En18 
    input [18:0] Wgt_8_360, // sfix19_En18 
    input [18:0] Wgt_8_361, // sfix19_En18 
    input [18:0] Wgt_8_362, // sfix19_En18 
    input [18:0] Wgt_8_363, // sfix19_En18 
    input [18:0] Wgt_8_364, // sfix19_En18 
    input [18:0] Wgt_8_365, // sfix19_En18 
    input [18:0] Wgt_8_366, // sfix19_En18 
    input [18:0] Wgt_8_367, // sfix19_En18 
    input [18:0] Wgt_8_368, // sfix19_En18 
    input [18:0] Wgt_8_369, // sfix19_En18 
    input [18:0] Wgt_8_370, // sfix19_En18 
    input [18:0] Wgt_8_371, // sfix19_En18 
    input [18:0] Wgt_8_372, // sfix19_En18 
    input [18:0] Wgt_8_373, // sfix19_En18 
    input [18:0] Wgt_8_374, // sfix19_En18 
    input [18:0] Wgt_8_375, // sfix19_En18 
    input [18:0] Wgt_8_376, // sfix19_En18 
    input [18:0] Wgt_8_377, // sfix19_En18 
    input [18:0] Wgt_8_378, // sfix19_En18 
    input [18:0] Wgt_8_379, // sfix19_En18 
    input [18:0] Wgt_8_380, // sfix19_En18 
    input [18:0] Wgt_8_381, // sfix19_En18 
    input [18:0] Wgt_8_382, // sfix19_En18 
    input [18:0] Wgt_8_383, // sfix19_En18 
    input [18:0] Wgt_8_384, // sfix19_En18 
    input [18:0] Wgt_8_385, // sfix19_En18 
    input [18:0] Wgt_8_386, // sfix19_En18 
    input [18:0] Wgt_8_387, // sfix19_En18 
    input [18:0] Wgt_8_388, // sfix19_En18 
    input [18:0] Wgt_8_389, // sfix19_En18 
    input [18:0] Wgt_8_390, // sfix19_En18 
    input [18:0] Wgt_8_391, // sfix19_En18 
    input [18:0] Wgt_8_392, // sfix19_En18 
    input [18:0] Wgt_8_393, // sfix19_En18 
    input [18:0] Wgt_8_394, // sfix19_En18 
    input [18:0] Wgt_8_395, // sfix19_En18 
    input [18:0] Wgt_8_396, // sfix19_En18 
    input [18:0] Wgt_8_397, // sfix19_En18 
    input [18:0] Wgt_8_398, // sfix19_En18 
    input [18:0] Wgt_8_399, // sfix19_En18 
    input [18:0] Wgt_8_400, // sfix19_En18 
    input [18:0] Wgt_8_401, // sfix19_En18 
    input [18:0] Wgt_8_402, // sfix19_En18 
    input [18:0] Wgt_8_403, // sfix19_En18 
    input [18:0] Wgt_8_404, // sfix19_En18 
    input [18:0] Wgt_8_405, // sfix19_En18 
    input [18:0] Wgt_8_406, // sfix19_En18 
    input [18:0] Wgt_8_407, // sfix19_En18 
    input [18:0] Wgt_8_408, // sfix19_En18 
    input [18:0] Wgt_8_409, // sfix19_En18 
    input [18:0] Wgt_8_410, // sfix19_En18 
    input [18:0] Wgt_8_411, // sfix19_En18 
    input [18:0] Wgt_8_412, // sfix19_En18 
    input [18:0] Wgt_8_413, // sfix19_En18 
    input [18:0] Wgt_8_414, // sfix19_En18 
    input [18:0] Wgt_8_415, // sfix19_En18 
    input [18:0] Wgt_8_416, // sfix19_En18 
    input [18:0] Wgt_8_417, // sfix19_En18 
    input [18:0] Wgt_8_418, // sfix19_En18 
    input [18:0] Wgt_8_419, // sfix19_En18 
    input [18:0] Wgt_8_420, // sfix19_En18 
    input [18:0] Wgt_8_421, // sfix19_En18 
    input [18:0] Wgt_8_422, // sfix19_En18 
    input [18:0] Wgt_8_423, // sfix19_En18 
    input [18:0] Wgt_8_424, // sfix19_En18 
    input [18:0] Wgt_8_425, // sfix19_En18 
    input [18:0] Wgt_8_426, // sfix19_En18 
    input [18:0] Wgt_8_427, // sfix19_En18 
    input [18:0] Wgt_8_428, // sfix19_En18 
    input [18:0] Wgt_8_429, // sfix19_En18 
    input [18:0] Wgt_8_430, // sfix19_En18 
    input [18:0] Wgt_8_431, // sfix19_En18 
    input [18:0] Wgt_8_432, // sfix19_En18 
    input [18:0] Wgt_8_433, // sfix19_En18 
    input [18:0] Wgt_8_434, // sfix19_En18 
    input [18:0] Wgt_8_435, // sfix19_En18 
    input [18:0] Wgt_8_436, // sfix19_En18 
    input [18:0] Wgt_8_437, // sfix19_En18 
    input [18:0] Wgt_8_438, // sfix19_En18 
    input [18:0] Wgt_8_439, // sfix19_En18 
    input [18:0] Wgt_8_440, // sfix19_En18 
    input [18:0] Wgt_8_441, // sfix19_En18 
    input [18:0] Wgt_8_442, // sfix19_En18 
    input [18:0] Wgt_8_443, // sfix19_En18 
    input [18:0] Wgt_8_444, // sfix19_En18 
    input [18:0] Wgt_8_445, // sfix19_En18 
    input [18:0] Wgt_8_446, // sfix19_En18 
    input [18:0] Wgt_8_447, // sfix19_En18 
    input [18:0] Wgt_8_448, // sfix19_En18 
    input [18:0] Wgt_8_449, // sfix19_En18 
    input [18:0] Wgt_8_450, // sfix19_En18 
    input [18:0] Wgt_8_451, // sfix19_En18 
    input [18:0] Wgt_8_452, // sfix19_En18 
    input [18:0] Wgt_8_453, // sfix19_En18 
    input [18:0] Wgt_8_454, // sfix19_En18 
    input [18:0] Wgt_8_455, // sfix19_En18 
    input [18:0] Wgt_8_456, // sfix19_En18 
    input [18:0] Wgt_8_457, // sfix19_En18 
    input [18:0] Wgt_8_458, // sfix19_En18 
    input [18:0] Wgt_8_459, // sfix19_En18 
    input [18:0] Wgt_8_460, // sfix19_En18 
    input [18:0] Wgt_8_461, // sfix19_En18 
    input [18:0] Wgt_8_462, // sfix19_En18 
    input [18:0] Wgt_8_463, // sfix19_En18 
    input [18:0] Wgt_8_464, // sfix19_En18 
    input [18:0] Wgt_8_465, // sfix19_En18 
    input [18:0] Wgt_8_466, // sfix19_En18 
    input [18:0] Wgt_8_467, // sfix19_En18 
    input [18:0] Wgt_8_468, // sfix19_En18 
    input [18:0] Wgt_8_469, // sfix19_En18 
    input [18:0] Wgt_8_470, // sfix19_En18 
    input [18:0] Wgt_8_471, // sfix19_En18 
    input [18:0] Wgt_8_472, // sfix19_En18 
    input [18:0] Wgt_8_473, // sfix19_En18 
    input [18:0] Wgt_8_474, // sfix19_En18 
    input [18:0] Wgt_8_475, // sfix19_En18 
    input [18:0] Wgt_8_476, // sfix19_En18 
    input [18:0] Wgt_8_477, // sfix19_En18 
    input [18:0] Wgt_8_478, // sfix19_En18 
    input [18:0] Wgt_8_479, // sfix19_En18 
    input [18:0] Wgt_8_480, // sfix19_En18 
    input [18:0] Wgt_8_481, // sfix19_En18 
    input [18:0] Wgt_8_482, // sfix19_En18 
    input [18:0] Wgt_8_483, // sfix19_En18 
    input [18:0] Wgt_8_484, // sfix19_En18 
    input [18:0] Wgt_8_485, // sfix19_En18 
    input [18:0] Wgt_8_486, // sfix19_En18 
    input [18:0] Wgt_8_487, // sfix19_En18 
    input [18:0] Wgt_8_488, // sfix19_En18 
    input [18:0] Wgt_8_489, // sfix19_En18 
    input [18:0] Wgt_8_490, // sfix19_En18 
    input [18:0] Wgt_8_491, // sfix19_En18 
    input [18:0] Wgt_8_492, // sfix19_En18 
    input [18:0] Wgt_8_493, // sfix19_En18 
    input [18:0] Wgt_8_494, // sfix19_En18 
    input [18:0] Wgt_8_495, // sfix19_En18 
    input [18:0] Wgt_8_496, // sfix19_En18 
    input [18:0] Wgt_8_497, // sfix19_En18 
    input [18:0] Wgt_8_498, // sfix19_En18 
    input [18:0] Wgt_8_499, // sfix19_En18 
    input [18:0] Wgt_8_500, // sfix19_En18 
    input [18:0] Wgt_8_501, // sfix19_En18 
    input [18:0] Wgt_8_502, // sfix19_En18 
    input [18:0] Wgt_8_503, // sfix19_En18 
    input [18:0] Wgt_8_504, // sfix19_En18 
    input [18:0] Wgt_8_505, // sfix19_En18 
    input [18:0] Wgt_8_506, // sfix19_En18 
    input [18:0] Wgt_8_507, // sfix19_En18 
    input [18:0] Wgt_8_508, // sfix19_En18 
    input [18:0] Wgt_8_509, // sfix19_En18 
    input [18:0] Wgt_8_510, // sfix19_En18 
    input [18:0] Wgt_8_511, // sfix19_En18 
    input [18:0] Wgt_8_512, // sfix19_En18 
    input [18:0] Wgt_8_513, // sfix19_En18 
    input [18:0] Wgt_8_514, // sfix19_En18 
    input [18:0] Wgt_8_515, // sfix19_En18 
    input [18:0] Wgt_8_516, // sfix19_En18 
    input [18:0] Wgt_8_517, // sfix19_En18 
    input [18:0] Wgt_8_518, // sfix19_En18 
    input [18:0] Wgt_8_519, // sfix19_En18 
    input [18:0] Wgt_8_520, // sfix19_En18 
    input [18:0] Wgt_8_521, // sfix19_En18 
    input [18:0] Wgt_8_522, // sfix19_En18 
    input [18:0] Wgt_8_523, // sfix19_En18 
    input [18:0] Wgt_8_524, // sfix19_En18 
    input [18:0] Wgt_8_525, // sfix19_En18 
    input [18:0] Wgt_8_526, // sfix19_En18 
    input [18:0] Wgt_8_527, // sfix19_En18 
    input [18:0] Wgt_8_528, // sfix19_En18 
    input [18:0] Wgt_8_529, // sfix19_En18 
    input [18:0] Wgt_8_530, // sfix19_En18 
    input [18:0] Wgt_8_531, // sfix19_En18 
    input [18:0] Wgt_8_532, // sfix19_En18 
    input [18:0] Wgt_8_533, // sfix19_En18 
    input [18:0] Wgt_8_534, // sfix19_En18 
    input [18:0] Wgt_8_535, // sfix19_En18 
    input [18:0] Wgt_8_536, // sfix19_En18 
    input [18:0] Wgt_8_537, // sfix19_En18 
    input [18:0] Wgt_8_538, // sfix19_En18 
    input [18:0] Wgt_8_539, // sfix19_En18 
    input [18:0] Wgt_8_540, // sfix19_En18 
    input [18:0] Wgt_8_541, // sfix19_En18 
    input [18:0] Wgt_8_542, // sfix19_En18 
    input [18:0] Wgt_8_543, // sfix19_En18 
    input [18:0] Wgt_8_544, // sfix19_En18 
    input [18:0] Wgt_8_545, // sfix19_En18 
    input [18:0] Wgt_8_546, // sfix19_En18 
    input [18:0] Wgt_8_547, // sfix19_En18 
    input [18:0] Wgt_8_548, // sfix19_En18 
    input [18:0] Wgt_8_549, // sfix19_En18 
    input [18:0] Wgt_8_550, // sfix19_En18 
    input [18:0] Wgt_8_551, // sfix19_En18 
    input [18:0] Wgt_8_552, // sfix19_En18 
    input [18:0] Wgt_8_553, // sfix19_En18 
    input [18:0] Wgt_8_554, // sfix19_En18 
    input [18:0] Wgt_8_555, // sfix19_En18 
    input [18:0] Wgt_8_556, // sfix19_En18 
    input [18:0] Wgt_8_557, // sfix19_En18 
    input [18:0] Wgt_8_558, // sfix19_En18 
    input [18:0] Wgt_8_559, // sfix19_En18 
    input [18:0] Wgt_8_560, // sfix19_En18 
    input [18:0] Wgt_8_561, // sfix19_En18 
    input [18:0] Wgt_8_562, // sfix19_En18 
    input [18:0] Wgt_8_563, // sfix19_En18 
    input [18:0] Wgt_8_564, // sfix19_En18 
    input [18:0] Wgt_8_565, // sfix19_En18 
    input [18:0] Wgt_8_566, // sfix19_En18 
    input [18:0] Wgt_8_567, // sfix19_En18 
    input [18:0] Wgt_8_568, // sfix19_En18 
    input [18:0] Wgt_8_569, // sfix19_En18 
    input [18:0] Wgt_8_570, // sfix19_En18 
    input [18:0] Wgt_8_571, // sfix19_En18 
    input [18:0] Wgt_8_572, // sfix19_En18 
    input [18:0] Wgt_8_573, // sfix19_En18 
    input [18:0] Wgt_8_574, // sfix19_En18 
    input [18:0] Wgt_8_575, // sfix19_En18 
    input [18:0] Wgt_8_576, // sfix19_En18 
    input [18:0] Wgt_8_577, // sfix19_En18 
    input [18:0] Wgt_8_578, // sfix19_En18 
    input [18:0] Wgt_8_579, // sfix19_En18 
    input [18:0] Wgt_8_580, // sfix19_En18 
    input [18:0] Wgt_8_581, // sfix19_En18 
    input [18:0] Wgt_8_582, // sfix19_En18 
    input [18:0] Wgt_8_583, // sfix19_En18 
    input [18:0] Wgt_8_584, // sfix19_En18 
    input [18:0] Wgt_8_585, // sfix19_En18 
    input [18:0] Wgt_8_586, // sfix19_En18 
    input [18:0] Wgt_8_587, // sfix19_En18 
    input [18:0] Wgt_8_588, // sfix19_En18 
    input [18:0] Wgt_8_589, // sfix19_En18 
    input [18:0] Wgt_8_590, // sfix19_En18 
    input [18:0] Wgt_8_591, // sfix19_En18 
    input [18:0] Wgt_8_592, // sfix19_En18 
    input [18:0] Wgt_8_593, // sfix19_En18 
    input [18:0] Wgt_8_594, // sfix19_En18 
    input [18:0] Wgt_8_595, // sfix19_En18 
    input [18:0] Wgt_8_596, // sfix19_En18 
    input [18:0] Wgt_8_597, // sfix19_En18 
    input [18:0] Wgt_8_598, // sfix19_En18 
    input [18:0] Wgt_8_599, // sfix19_En18 
    input [18:0] Wgt_8_600, // sfix19_En18 
    input [18:0] Wgt_8_601, // sfix19_En18 
    input [18:0] Wgt_8_602, // sfix19_En18 
    input [18:0] Wgt_8_603, // sfix19_En18 
    input [18:0] Wgt_8_604, // sfix19_En18 
    input [18:0] Wgt_8_605, // sfix19_En18 
    input [18:0] Wgt_8_606, // sfix19_En18 
    input [18:0] Wgt_8_607, // sfix19_En18 
    input [18:0] Wgt_8_608, // sfix19_En18 
    input [18:0] Wgt_8_609, // sfix19_En18 
    input [18:0] Wgt_8_610, // sfix19_En18 
    input [18:0] Wgt_8_611, // sfix19_En18 
    input [18:0] Wgt_8_612, // sfix19_En18 
    input [18:0] Wgt_8_613, // sfix19_En18 
    input [18:0] Wgt_8_614, // sfix19_En18 
    input [18:0] Wgt_8_615, // sfix19_En18 
    input [18:0] Wgt_8_616, // sfix19_En18 
    input [18:0] Wgt_8_617, // sfix19_En18 
    input [18:0] Wgt_8_618, // sfix19_En18 
    input [18:0] Wgt_8_619, // sfix19_En18 
    input [18:0] Wgt_8_620, // sfix19_En18 
    input [18:0] Wgt_8_621, // sfix19_En18 
    input [18:0] Wgt_8_622, // sfix19_En18 
    input [18:0] Wgt_8_623, // sfix19_En18 
    input [18:0] Wgt_8_624, // sfix19_En18 
    input [18:0] Wgt_8_625, // sfix19_En18 
    input [18:0] Wgt_8_626, // sfix19_En18 
    input [18:0] Wgt_8_627, // sfix19_En18 
    input [18:0] Wgt_8_628, // sfix19_En18 
    input [18:0] Wgt_8_629, // sfix19_En18 
    input [18:0] Wgt_8_630, // sfix19_En18 
    input [18:0] Wgt_8_631, // sfix19_En18 
    input [18:0] Wgt_8_632, // sfix19_En18 
    input [18:0] Wgt_8_633, // sfix19_En18 
    input [18:0] Wgt_8_634, // sfix19_En18 
    input [18:0] Wgt_8_635, // sfix19_En18 
    input [18:0] Wgt_8_636, // sfix19_En18 
    input [18:0] Wgt_8_637, // sfix19_En18 
    input [18:0] Wgt_8_638, // sfix19_En18 
    input [18:0] Wgt_8_639, // sfix19_En18 
    input [18:0] Wgt_8_640, // sfix19_En18 
    input [18:0] Wgt_8_641, // sfix19_En18 
    input [18:0] Wgt_8_642, // sfix19_En18 
    input [18:0] Wgt_8_643, // sfix19_En18 
    input [18:0] Wgt_8_644, // sfix19_En18 
    input [18:0] Wgt_8_645, // sfix19_En18 
    input [18:0] Wgt_8_646, // sfix19_En18 
    input [18:0] Wgt_8_647, // sfix19_En18 
    input [18:0] Wgt_8_648, // sfix19_En18 
    input [18:0] Wgt_8_649, // sfix19_En18 
    input [18:0] Wgt_8_650, // sfix19_En18 
    input [18:0] Wgt_8_651, // sfix19_En18 
    input [18:0] Wgt_8_652, // sfix19_En18 
    input [18:0] Wgt_8_653, // sfix19_En18 
    input [18:0] Wgt_8_654, // sfix19_En18 
    input [18:0] Wgt_8_655, // sfix19_En18 
    input [18:0] Wgt_8_656, // sfix19_En18 
    input [18:0] Wgt_8_657, // sfix19_En18 
    input [18:0] Wgt_8_658, // sfix19_En18 
    input [18:0] Wgt_8_659, // sfix19_En18 
    input [18:0] Wgt_8_660, // sfix19_En18 
    input [18:0] Wgt_8_661, // sfix19_En18 
    input [18:0] Wgt_8_662, // sfix19_En18 
    input [18:0] Wgt_8_663, // sfix19_En18 
    input [18:0] Wgt_8_664, // sfix19_En18 
    input [18:0] Wgt_8_665, // sfix19_En18 
    input [18:0] Wgt_8_666, // sfix19_En18 
    input [18:0] Wgt_8_667, // sfix19_En18 
    input [18:0] Wgt_8_668, // sfix19_En18 
    input [18:0] Wgt_8_669, // sfix19_En18 
    input [18:0] Wgt_8_670, // sfix19_En18 
    input [18:0] Wgt_8_671, // sfix19_En18 
    input [18:0] Wgt_8_672, // sfix19_En18 
    input [18:0] Wgt_8_673, // sfix19_En18 
    input [18:0] Wgt_8_674, // sfix19_En18 
    input [18:0] Wgt_8_675, // sfix19_En18 
    input [18:0] Wgt_8_676, // sfix19_En18 
    input [18:0] Wgt_8_677, // sfix19_En18 
    input [18:0] Wgt_8_678, // sfix19_En18 
    input [18:0] Wgt_8_679, // sfix19_En18 
    input [18:0] Wgt_8_680, // sfix19_En18 
    input [18:0] Wgt_8_681, // sfix19_En18 
    input [18:0] Wgt_8_682, // sfix19_En18 
    input [18:0] Wgt_8_683, // sfix19_En18 
    input [18:0] Wgt_8_684, // sfix19_En18 
    input [18:0] Wgt_8_685, // sfix19_En18 
    input [18:0] Wgt_8_686, // sfix19_En18 
    input [18:0] Wgt_8_687, // sfix19_En18 
    input [18:0] Wgt_8_688, // sfix19_En18 
    input [18:0] Wgt_8_689, // sfix19_En18 
    input [18:0] Wgt_8_690, // sfix19_En18 
    input [18:0] Wgt_8_691, // sfix19_En18 
    input [18:0] Wgt_8_692, // sfix19_En18 
    input [18:0] Wgt_8_693, // sfix19_En18 
    input [18:0] Wgt_8_694, // sfix19_En18 
    input [18:0] Wgt_8_695, // sfix19_En18 
    input [18:0] Wgt_8_696, // sfix19_En18 
    input [18:0] Wgt_8_697, // sfix19_En18 
    input [18:0] Wgt_8_698, // sfix19_En18 
    input [18:0] Wgt_8_699, // sfix19_En18 
    input [18:0] Wgt_8_700, // sfix19_En18 
    input [18:0] Wgt_8_701, // sfix19_En18 
    input [18:0] Wgt_8_702, // sfix19_En18 
    input [18:0] Wgt_8_703, // sfix19_En18 
    input [18:0] Wgt_8_704, // sfix19_En18 
    input [18:0] Wgt_8_705, // sfix19_En18 
    input [18:0] Wgt_8_706, // sfix19_En18 
    input [18:0] Wgt_8_707, // sfix19_En18 
    input [18:0] Wgt_8_708, // sfix19_En18 
    input [18:0] Wgt_8_709, // sfix19_En18 
    input [18:0] Wgt_8_710, // sfix19_En18 
    input [18:0] Wgt_8_711, // sfix19_En18 
    input [18:0] Wgt_8_712, // sfix19_En18 
    input [18:0] Wgt_8_713, // sfix19_En18 
    input [18:0] Wgt_8_714, // sfix19_En18 
    input [18:0] Wgt_8_715, // sfix19_En18 
    input [18:0] Wgt_8_716, // sfix19_En18 
    input [18:0] Wgt_8_717, // sfix19_En18 
    input [18:0] Wgt_8_718, // sfix19_En18 
    input [18:0] Wgt_8_719, // sfix19_En18 
    input [18:0] Wgt_8_720, // sfix19_En18 
    input [18:0] Wgt_8_721, // sfix19_En18 
    input [18:0] Wgt_8_722, // sfix19_En18 
    input [18:0] Wgt_8_723, // sfix19_En18 
    input [18:0] Wgt_8_724, // sfix19_En18 
    input [18:0] Wgt_8_725, // sfix19_En18 
    input [18:0] Wgt_8_726, // sfix19_En18 
    input [18:0] Wgt_8_727, // sfix19_En18 
    input [18:0] Wgt_8_728, // sfix19_En18 
    input [18:0] Wgt_8_729, // sfix19_En18 
    input [18:0] Wgt_8_730, // sfix19_En18 
    input [18:0] Wgt_8_731, // sfix19_En18 
    input [18:0] Wgt_8_732, // sfix19_En18 
    input [18:0] Wgt_8_733, // sfix19_En18 
    input [18:0] Wgt_8_734, // sfix19_En18 
    input [18:0] Wgt_8_735, // sfix19_En18 
    input [18:0] Wgt_8_736, // sfix19_En18 
    input [18:0] Wgt_8_737, // sfix19_En18 
    input [18:0] Wgt_8_738, // sfix19_En18 
    input [18:0] Wgt_8_739, // sfix19_En18 
    input [18:0] Wgt_8_740, // sfix19_En18 
    input [18:0] Wgt_8_741, // sfix19_En18 
    input [18:0] Wgt_8_742, // sfix19_En18 
    input [18:0] Wgt_8_743, // sfix19_En18 
    input [18:0] Wgt_8_744, // sfix19_En18 
    input [18:0] Wgt_8_745, // sfix19_En18 
    input [18:0] Wgt_8_746, // sfix19_En18 
    input [18:0] Wgt_8_747, // sfix19_En18 
    input [18:0] Wgt_8_748, // sfix19_En18 
    input [18:0] Wgt_8_749, // sfix19_En18 
    input [18:0] Wgt_8_750, // sfix19_En18 
    input [18:0] Wgt_8_751, // sfix19_En18 
    input [18:0] Wgt_8_752, // sfix19_En18 
    input [18:0] Wgt_8_753, // sfix19_En18 
    input [18:0] Wgt_8_754, // sfix19_En18 
    input [18:0] Wgt_8_755, // sfix19_En18 
    input [18:0] Wgt_8_756, // sfix19_En18 
    input [18:0] Wgt_8_757, // sfix19_En18 
    input [18:0] Wgt_8_758, // sfix19_En18 
    input [18:0] Wgt_8_759, // sfix19_En18 
    input [18:0] Wgt_8_760, // sfix19_En18 
    input [18:0] Wgt_8_761, // sfix19_En18 
    input [18:0] Wgt_8_762, // sfix19_En18 
    input [18:0] Wgt_8_763, // sfix19_En18 
    input [18:0] Wgt_8_764, // sfix19_En18 
    input [18:0] Wgt_8_765, // sfix19_En18 
    input [18:0] Wgt_8_766, // sfix19_En18 
    input [18:0] Wgt_8_767, // sfix19_En18 
    input [18:0] Wgt_8_768, // sfix19_En18 
    input [18:0] Wgt_8_769, // sfix19_En18 
    input [18:0] Wgt_8_770, // sfix19_En18 
    input [18:0] Wgt_8_771, // sfix19_En18 
    input [18:0] Wgt_8_772, // sfix19_En18 
    input [18:0] Wgt_8_773, // sfix19_En18 
    input [18:0] Wgt_8_774, // sfix19_En18 
    input [18:0] Wgt_8_775, // sfix19_En18 
    input [18:0] Wgt_8_776, // sfix19_En18 
    input [18:0] Wgt_8_777, // sfix19_En18 
    input [18:0] Wgt_8_778, // sfix19_En18 
    input [18:0] Wgt_8_779, // sfix19_En18 
    input [18:0] Wgt_8_780, // sfix19_En18 
    input [18:0] Wgt_8_781, // sfix19_En18 
    input [18:0] Wgt_8_782, // sfix19_En18 
    input [18:0] Wgt_8_783, // sfix19_En18 
    input [18:0] Wgt_8_784, // sfix19_En18 
    input [18:0] Wgt_9_0, // sfix19_En18 
    input [18:0] Wgt_9_1, // sfix19_En18 
    input [18:0] Wgt_9_2, // sfix19_En18 
    input [18:0] Wgt_9_3, // sfix19_En18 
    input [18:0] Wgt_9_4, // sfix19_En18 
    input [18:0] Wgt_9_5, // sfix19_En18 
    input [18:0] Wgt_9_6, // sfix19_En18 
    input [18:0] Wgt_9_7, // sfix19_En18 
    input [18:0] Wgt_9_8, // sfix19_En18 
    input [18:0] Wgt_9_9, // sfix19_En18 
    input [18:0] Wgt_9_10, // sfix19_En18 
    input [18:0] Wgt_9_11, // sfix19_En18 
    input [18:0] Wgt_9_12, // sfix19_En18 
    input [18:0] Wgt_9_13, // sfix19_En18 
    input [18:0] Wgt_9_14, // sfix19_En18 
    input [18:0] Wgt_9_15, // sfix19_En18 
    input [18:0] Wgt_9_16, // sfix19_En18 
    input [18:0] Wgt_9_17, // sfix19_En18 
    input [18:0] Wgt_9_18, // sfix19_En18 
    input [18:0] Wgt_9_19, // sfix19_En18 
    input [18:0] Wgt_9_20, // sfix19_En18 
    input [18:0] Wgt_9_21, // sfix19_En18 
    input [18:0] Wgt_9_22, // sfix19_En18 
    input [18:0] Wgt_9_23, // sfix19_En18 
    input [18:0] Wgt_9_24, // sfix19_En18 
    input [18:0] Wgt_9_25, // sfix19_En18 
    input [18:0] Wgt_9_26, // sfix19_En18 
    input [18:0] Wgt_9_27, // sfix19_En18 
    input [18:0] Wgt_9_28, // sfix19_En18 
    input [18:0] Wgt_9_29, // sfix19_En18 
    input [18:0] Wgt_9_30, // sfix19_En18 
    input [18:0] Wgt_9_31, // sfix19_En18 
    input [18:0] Wgt_9_32, // sfix19_En18 
    input [18:0] Wgt_9_33, // sfix19_En18 
    input [18:0] Wgt_9_34, // sfix19_En18 
    input [18:0] Wgt_9_35, // sfix19_En18 
    input [18:0] Wgt_9_36, // sfix19_En18 
    input [18:0] Wgt_9_37, // sfix19_En18 
    input [18:0] Wgt_9_38, // sfix19_En18 
    input [18:0] Wgt_9_39, // sfix19_En18 
    input [18:0] Wgt_9_40, // sfix19_En18 
    input [18:0] Wgt_9_41, // sfix19_En18 
    input [18:0] Wgt_9_42, // sfix19_En18 
    input [18:0] Wgt_9_43, // sfix19_En18 
    input [18:0] Wgt_9_44, // sfix19_En18 
    input [18:0] Wgt_9_45, // sfix19_En18 
    input [18:0] Wgt_9_46, // sfix19_En18 
    input [18:0] Wgt_9_47, // sfix19_En18 
    input [18:0] Wgt_9_48, // sfix19_En18 
    input [18:0] Wgt_9_49, // sfix19_En18 
    input [18:0] Wgt_9_50, // sfix19_En18 
    input [18:0] Wgt_9_51, // sfix19_En18 
    input [18:0] Wgt_9_52, // sfix19_En18 
    input [18:0] Wgt_9_53, // sfix19_En18 
    input [18:0] Wgt_9_54, // sfix19_En18 
    input [18:0] Wgt_9_55, // sfix19_En18 
    input [18:0] Wgt_9_56, // sfix19_En18 
    input [18:0] Wgt_9_57, // sfix19_En18 
    input [18:0] Wgt_9_58, // sfix19_En18 
    input [18:0] Wgt_9_59, // sfix19_En18 
    input [18:0] Wgt_9_60, // sfix19_En18 
    input [18:0] Wgt_9_61, // sfix19_En18 
    input [18:0] Wgt_9_62, // sfix19_En18 
    input [18:0] Wgt_9_63, // sfix19_En18 
    input [18:0] Wgt_9_64, // sfix19_En18 
    input [18:0] Wgt_9_65, // sfix19_En18 
    input [18:0] Wgt_9_66, // sfix19_En18 
    input [18:0] Wgt_9_67, // sfix19_En18 
    input [18:0] Wgt_9_68, // sfix19_En18 
    input [18:0] Wgt_9_69, // sfix19_En18 
    input [18:0] Wgt_9_70, // sfix19_En18 
    input [18:0] Wgt_9_71, // sfix19_En18 
    input [18:0] Wgt_9_72, // sfix19_En18 
    input [18:0] Wgt_9_73, // sfix19_En18 
    input [18:0] Wgt_9_74, // sfix19_En18 
    input [18:0] Wgt_9_75, // sfix19_En18 
    input [18:0] Wgt_9_76, // sfix19_En18 
    input [18:0] Wgt_9_77, // sfix19_En18 
    input [18:0] Wgt_9_78, // sfix19_En18 
    input [18:0] Wgt_9_79, // sfix19_En18 
    input [18:0] Wgt_9_80, // sfix19_En18 
    input [18:0] Wgt_9_81, // sfix19_En18 
    input [18:0] Wgt_9_82, // sfix19_En18 
    input [18:0] Wgt_9_83, // sfix19_En18 
    input [18:0] Wgt_9_84, // sfix19_En18 
    input [18:0] Wgt_9_85, // sfix19_En18 
    input [18:0] Wgt_9_86, // sfix19_En18 
    input [18:0] Wgt_9_87, // sfix19_En18 
    input [18:0] Wgt_9_88, // sfix19_En18 
    input [18:0] Wgt_9_89, // sfix19_En18 
    input [18:0] Wgt_9_90, // sfix19_En18 
    input [18:0] Wgt_9_91, // sfix19_En18 
    input [18:0] Wgt_9_92, // sfix19_En18 
    input [18:0] Wgt_9_93, // sfix19_En18 
    input [18:0] Wgt_9_94, // sfix19_En18 
    input [18:0] Wgt_9_95, // sfix19_En18 
    input [18:0] Wgt_9_96, // sfix19_En18 
    input [18:0] Wgt_9_97, // sfix19_En18 
    input [18:0] Wgt_9_98, // sfix19_En18 
    input [18:0] Wgt_9_99, // sfix19_En18 
    input [18:0] Wgt_9_100, // sfix19_En18 
    input [18:0] Wgt_9_101, // sfix19_En18 
    input [18:0] Wgt_9_102, // sfix19_En18 
    input [18:0] Wgt_9_103, // sfix19_En18 
    input [18:0] Wgt_9_104, // sfix19_En18 
    input [18:0] Wgt_9_105, // sfix19_En18 
    input [18:0] Wgt_9_106, // sfix19_En18 
    input [18:0] Wgt_9_107, // sfix19_En18 
    input [18:0] Wgt_9_108, // sfix19_En18 
    input [18:0] Wgt_9_109, // sfix19_En18 
    input [18:0] Wgt_9_110, // sfix19_En18 
    input [18:0] Wgt_9_111, // sfix19_En18 
    input [18:0] Wgt_9_112, // sfix19_En18 
    input [18:0] Wgt_9_113, // sfix19_En18 
    input [18:0] Wgt_9_114, // sfix19_En18 
    input [18:0] Wgt_9_115, // sfix19_En18 
    input [18:0] Wgt_9_116, // sfix19_En18 
    input [18:0] Wgt_9_117, // sfix19_En18 
    input [18:0] Wgt_9_118, // sfix19_En18 
    input [18:0] Wgt_9_119, // sfix19_En18 
    input [18:0] Wgt_9_120, // sfix19_En18 
    input [18:0] Wgt_9_121, // sfix19_En18 
    input [18:0] Wgt_9_122, // sfix19_En18 
    input [18:0] Wgt_9_123, // sfix19_En18 
    input [18:0] Wgt_9_124, // sfix19_En18 
    input [18:0] Wgt_9_125, // sfix19_En18 
    input [18:0] Wgt_9_126, // sfix19_En18 
    input [18:0] Wgt_9_127, // sfix19_En18 
    input [18:0] Wgt_9_128, // sfix19_En18 
    input [18:0] Wgt_9_129, // sfix19_En18 
    input [18:0] Wgt_9_130, // sfix19_En18 
    input [18:0] Wgt_9_131, // sfix19_En18 
    input [18:0] Wgt_9_132, // sfix19_En18 
    input [18:0] Wgt_9_133, // sfix19_En18 
    input [18:0] Wgt_9_134, // sfix19_En18 
    input [18:0] Wgt_9_135, // sfix19_En18 
    input [18:0] Wgt_9_136, // sfix19_En18 
    input [18:0] Wgt_9_137, // sfix19_En18 
    input [18:0] Wgt_9_138, // sfix19_En18 
    input [18:0] Wgt_9_139, // sfix19_En18 
    input [18:0] Wgt_9_140, // sfix19_En18 
    input [18:0] Wgt_9_141, // sfix19_En18 
    input [18:0] Wgt_9_142, // sfix19_En18 
    input [18:0] Wgt_9_143, // sfix19_En18 
    input [18:0] Wgt_9_144, // sfix19_En18 
    input [18:0] Wgt_9_145, // sfix19_En18 
    input [18:0] Wgt_9_146, // sfix19_En18 
    input [18:0] Wgt_9_147, // sfix19_En18 
    input [18:0] Wgt_9_148, // sfix19_En18 
    input [18:0] Wgt_9_149, // sfix19_En18 
    input [18:0] Wgt_9_150, // sfix19_En18 
    input [18:0] Wgt_9_151, // sfix19_En18 
    input [18:0] Wgt_9_152, // sfix19_En18 
    input [18:0] Wgt_9_153, // sfix19_En18 
    input [18:0] Wgt_9_154, // sfix19_En18 
    input [18:0] Wgt_9_155, // sfix19_En18 
    input [18:0] Wgt_9_156, // sfix19_En18 
    input [18:0] Wgt_9_157, // sfix19_En18 
    input [18:0] Wgt_9_158, // sfix19_En18 
    input [18:0] Wgt_9_159, // sfix19_En18 
    input [18:0] Wgt_9_160, // sfix19_En18 
    input [18:0] Wgt_9_161, // sfix19_En18 
    input [18:0] Wgt_9_162, // sfix19_En18 
    input [18:0] Wgt_9_163, // sfix19_En18 
    input [18:0] Wgt_9_164, // sfix19_En18 
    input [18:0] Wgt_9_165, // sfix19_En18 
    input [18:0] Wgt_9_166, // sfix19_En18 
    input [18:0] Wgt_9_167, // sfix19_En18 
    input [18:0] Wgt_9_168, // sfix19_En18 
    input [18:0] Wgt_9_169, // sfix19_En18 
    input [18:0] Wgt_9_170, // sfix19_En18 
    input [18:0] Wgt_9_171, // sfix19_En18 
    input [18:0] Wgt_9_172, // sfix19_En18 
    input [18:0] Wgt_9_173, // sfix19_En18 
    input [18:0] Wgt_9_174, // sfix19_En18 
    input [18:0] Wgt_9_175, // sfix19_En18 
    input [18:0] Wgt_9_176, // sfix19_En18 
    input [18:0] Wgt_9_177, // sfix19_En18 
    input [18:0] Wgt_9_178, // sfix19_En18 
    input [18:0] Wgt_9_179, // sfix19_En18 
    input [18:0] Wgt_9_180, // sfix19_En18 
    input [18:0] Wgt_9_181, // sfix19_En18 
    input [18:0] Wgt_9_182, // sfix19_En18 
    input [18:0] Wgt_9_183, // sfix19_En18 
    input [18:0] Wgt_9_184, // sfix19_En18 
    input [18:0] Wgt_9_185, // sfix19_En18 
    input [18:0] Wgt_9_186, // sfix19_En18 
    input [18:0] Wgt_9_187, // sfix19_En18 
    input [18:0] Wgt_9_188, // sfix19_En18 
    input [18:0] Wgt_9_189, // sfix19_En18 
    input [18:0] Wgt_9_190, // sfix19_En18 
    input [18:0] Wgt_9_191, // sfix19_En18 
    input [18:0] Wgt_9_192, // sfix19_En18 
    input [18:0] Wgt_9_193, // sfix19_En18 
    input [18:0] Wgt_9_194, // sfix19_En18 
    input [18:0] Wgt_9_195, // sfix19_En18 
    input [18:0] Wgt_9_196, // sfix19_En18 
    input [18:0] Wgt_9_197, // sfix19_En18 
    input [18:0] Wgt_9_198, // sfix19_En18 
    input [18:0] Wgt_9_199, // sfix19_En18 
    input [18:0] Wgt_9_200, // sfix19_En18 
    input [18:0] Wgt_9_201, // sfix19_En18 
    input [18:0] Wgt_9_202, // sfix19_En18 
    input [18:0] Wgt_9_203, // sfix19_En18 
    input [18:0] Wgt_9_204, // sfix19_En18 
    input [18:0] Wgt_9_205, // sfix19_En18 
    input [18:0] Wgt_9_206, // sfix19_En18 
    input [18:0] Wgt_9_207, // sfix19_En18 
    input [18:0] Wgt_9_208, // sfix19_En18 
    input [18:0] Wgt_9_209, // sfix19_En18 
    input [18:0] Wgt_9_210, // sfix19_En18 
    input [18:0] Wgt_9_211, // sfix19_En18 
    input [18:0] Wgt_9_212, // sfix19_En18 
    input [18:0] Wgt_9_213, // sfix19_En18 
    input [18:0] Wgt_9_214, // sfix19_En18 
    input [18:0] Wgt_9_215, // sfix19_En18 
    input [18:0] Wgt_9_216, // sfix19_En18 
    input [18:0] Wgt_9_217, // sfix19_En18 
    input [18:0] Wgt_9_218, // sfix19_En18 
    input [18:0] Wgt_9_219, // sfix19_En18 
    input [18:0] Wgt_9_220, // sfix19_En18 
    input [18:0] Wgt_9_221, // sfix19_En18 
    input [18:0] Wgt_9_222, // sfix19_En18 
    input [18:0] Wgt_9_223, // sfix19_En18 
    input [18:0] Wgt_9_224, // sfix19_En18 
    input [18:0] Wgt_9_225, // sfix19_En18 
    input [18:0] Wgt_9_226, // sfix19_En18 
    input [18:0] Wgt_9_227, // sfix19_En18 
    input [18:0] Wgt_9_228, // sfix19_En18 
    input [18:0] Wgt_9_229, // sfix19_En18 
    input [18:0] Wgt_9_230, // sfix19_En18 
    input [18:0] Wgt_9_231, // sfix19_En18 
    input [18:0] Wgt_9_232, // sfix19_En18 
    input [18:0] Wgt_9_233, // sfix19_En18 
    input [18:0] Wgt_9_234, // sfix19_En18 
    input [18:0] Wgt_9_235, // sfix19_En18 
    input [18:0] Wgt_9_236, // sfix19_En18 
    input [18:0] Wgt_9_237, // sfix19_En18 
    input [18:0] Wgt_9_238, // sfix19_En18 
    input [18:0] Wgt_9_239, // sfix19_En18 
    input [18:0] Wgt_9_240, // sfix19_En18 
    input [18:0] Wgt_9_241, // sfix19_En18 
    input [18:0] Wgt_9_242, // sfix19_En18 
    input [18:0] Wgt_9_243, // sfix19_En18 
    input [18:0] Wgt_9_244, // sfix19_En18 
    input [18:0] Wgt_9_245, // sfix19_En18 
    input [18:0] Wgt_9_246, // sfix19_En18 
    input [18:0] Wgt_9_247, // sfix19_En18 
    input [18:0] Wgt_9_248, // sfix19_En18 
    input [18:0] Wgt_9_249, // sfix19_En18 
    input [18:0] Wgt_9_250, // sfix19_En18 
    input [18:0] Wgt_9_251, // sfix19_En18 
    input [18:0] Wgt_9_252, // sfix19_En18 
    input [18:0] Wgt_9_253, // sfix19_En18 
    input [18:0] Wgt_9_254, // sfix19_En18 
    input [18:0] Wgt_9_255, // sfix19_En18 
    input [18:0] Wgt_9_256, // sfix19_En18 
    input [18:0] Wgt_9_257, // sfix19_En18 
    input [18:0] Wgt_9_258, // sfix19_En18 
    input [18:0] Wgt_9_259, // sfix19_En18 
    input [18:0] Wgt_9_260, // sfix19_En18 
    input [18:0] Wgt_9_261, // sfix19_En18 
    input [18:0] Wgt_9_262, // sfix19_En18 
    input [18:0] Wgt_9_263, // sfix19_En18 
    input [18:0] Wgt_9_264, // sfix19_En18 
    input [18:0] Wgt_9_265, // sfix19_En18 
    input [18:0] Wgt_9_266, // sfix19_En18 
    input [18:0] Wgt_9_267, // sfix19_En18 
    input [18:0] Wgt_9_268, // sfix19_En18 
    input [18:0] Wgt_9_269, // sfix19_En18 
    input [18:0] Wgt_9_270, // sfix19_En18 
    input [18:0] Wgt_9_271, // sfix19_En18 
    input [18:0] Wgt_9_272, // sfix19_En18 
    input [18:0] Wgt_9_273, // sfix19_En18 
    input [18:0] Wgt_9_274, // sfix19_En18 
    input [18:0] Wgt_9_275, // sfix19_En18 
    input [18:0] Wgt_9_276, // sfix19_En18 
    input [18:0] Wgt_9_277, // sfix19_En18 
    input [18:0] Wgt_9_278, // sfix19_En18 
    input [18:0] Wgt_9_279, // sfix19_En18 
    input [18:0] Wgt_9_280, // sfix19_En18 
    input [18:0] Wgt_9_281, // sfix19_En18 
    input [18:0] Wgt_9_282, // sfix19_En18 
    input [18:0] Wgt_9_283, // sfix19_En18 
    input [18:0] Wgt_9_284, // sfix19_En18 
    input [18:0] Wgt_9_285, // sfix19_En18 
    input [18:0] Wgt_9_286, // sfix19_En18 
    input [18:0] Wgt_9_287, // sfix19_En18 
    input [18:0] Wgt_9_288, // sfix19_En18 
    input [18:0] Wgt_9_289, // sfix19_En18 
    input [18:0] Wgt_9_290, // sfix19_En18 
    input [18:0] Wgt_9_291, // sfix19_En18 
    input [18:0] Wgt_9_292, // sfix19_En18 
    input [18:0] Wgt_9_293, // sfix19_En18 
    input [18:0] Wgt_9_294, // sfix19_En18 
    input [18:0] Wgt_9_295, // sfix19_En18 
    input [18:0] Wgt_9_296, // sfix19_En18 
    input [18:0] Wgt_9_297, // sfix19_En18 
    input [18:0] Wgt_9_298, // sfix19_En18 
    input [18:0] Wgt_9_299, // sfix19_En18 
    input [18:0] Wgt_9_300, // sfix19_En18 
    input [18:0] Wgt_9_301, // sfix19_En18 
    input [18:0] Wgt_9_302, // sfix19_En18 
    input [18:0] Wgt_9_303, // sfix19_En18 
    input [18:0] Wgt_9_304, // sfix19_En18 
    input [18:0] Wgt_9_305, // sfix19_En18 
    input [18:0] Wgt_9_306, // sfix19_En18 
    input [18:0] Wgt_9_307, // sfix19_En18 
    input [18:0] Wgt_9_308, // sfix19_En18 
    input [18:0] Wgt_9_309, // sfix19_En18 
    input [18:0] Wgt_9_310, // sfix19_En18 
    input [18:0] Wgt_9_311, // sfix19_En18 
    input [18:0] Wgt_9_312, // sfix19_En18 
    input [18:0] Wgt_9_313, // sfix19_En18 
    input [18:0] Wgt_9_314, // sfix19_En18 
    input [18:0] Wgt_9_315, // sfix19_En18 
    input [18:0] Wgt_9_316, // sfix19_En18 
    input [18:0] Wgt_9_317, // sfix19_En18 
    input [18:0] Wgt_9_318, // sfix19_En18 
    input [18:0] Wgt_9_319, // sfix19_En18 
    input [18:0] Wgt_9_320, // sfix19_En18 
    input [18:0] Wgt_9_321, // sfix19_En18 
    input [18:0] Wgt_9_322, // sfix19_En18 
    input [18:0] Wgt_9_323, // sfix19_En18 
    input [18:0] Wgt_9_324, // sfix19_En18 
    input [18:0] Wgt_9_325, // sfix19_En18 
    input [18:0] Wgt_9_326, // sfix19_En18 
    input [18:0] Wgt_9_327, // sfix19_En18 
    input [18:0] Wgt_9_328, // sfix19_En18 
    input [18:0] Wgt_9_329, // sfix19_En18 
    input [18:0] Wgt_9_330, // sfix19_En18 
    input [18:0] Wgt_9_331, // sfix19_En18 
    input [18:0] Wgt_9_332, // sfix19_En18 
    input [18:0] Wgt_9_333, // sfix19_En18 
    input [18:0] Wgt_9_334, // sfix19_En18 
    input [18:0] Wgt_9_335, // sfix19_En18 
    input [18:0] Wgt_9_336, // sfix19_En18 
    input [18:0] Wgt_9_337, // sfix19_En18 
    input [18:0] Wgt_9_338, // sfix19_En18 
    input [18:0] Wgt_9_339, // sfix19_En18 
    input [18:0] Wgt_9_340, // sfix19_En18 
    input [18:0] Wgt_9_341, // sfix19_En18 
    input [18:0] Wgt_9_342, // sfix19_En18 
    input [18:0] Wgt_9_343, // sfix19_En18 
    input [18:0] Wgt_9_344, // sfix19_En18 
    input [18:0] Wgt_9_345, // sfix19_En18 
    input [18:0] Wgt_9_346, // sfix19_En18 
    input [18:0] Wgt_9_347, // sfix19_En18 
    input [18:0] Wgt_9_348, // sfix19_En18 
    input [18:0] Wgt_9_349, // sfix19_En18 
    input [18:0] Wgt_9_350, // sfix19_En18 
    input [18:0] Wgt_9_351, // sfix19_En18 
    input [18:0] Wgt_9_352, // sfix19_En18 
    input [18:0] Wgt_9_353, // sfix19_En18 
    input [18:0] Wgt_9_354, // sfix19_En18 
    input [18:0] Wgt_9_355, // sfix19_En18 
    input [18:0] Wgt_9_356, // sfix19_En18 
    input [18:0] Wgt_9_357, // sfix19_En18 
    input [18:0] Wgt_9_358, // sfix19_En18 
    input [18:0] Wgt_9_359, // sfix19_En18 
    input [18:0] Wgt_9_360, // sfix19_En18 
    input [18:0] Wgt_9_361, // sfix19_En18 
    input [18:0] Wgt_9_362, // sfix19_En18 
    input [18:0] Wgt_9_363, // sfix19_En18 
    input [18:0] Wgt_9_364, // sfix19_En18 
    input [18:0] Wgt_9_365, // sfix19_En18 
    input [18:0] Wgt_9_366, // sfix19_En18 
    input [18:0] Wgt_9_367, // sfix19_En18 
    input [18:0] Wgt_9_368, // sfix19_En18 
    input [18:0] Wgt_9_369, // sfix19_En18 
    input [18:0] Wgt_9_370, // sfix19_En18 
    input [18:0] Wgt_9_371, // sfix19_En18 
    input [18:0] Wgt_9_372, // sfix19_En18 
    input [18:0] Wgt_9_373, // sfix19_En18 
    input [18:0] Wgt_9_374, // sfix19_En18 
    input [18:0] Wgt_9_375, // sfix19_En18 
    input [18:0] Wgt_9_376, // sfix19_En18 
    input [18:0] Wgt_9_377, // sfix19_En18 
    input [18:0] Wgt_9_378, // sfix19_En18 
    input [18:0] Wgt_9_379, // sfix19_En18 
    input [18:0] Wgt_9_380, // sfix19_En18 
    input [18:0] Wgt_9_381, // sfix19_En18 
    input [18:0] Wgt_9_382, // sfix19_En18 
    input [18:0] Wgt_9_383, // sfix19_En18 
    input [18:0] Wgt_9_384, // sfix19_En18 
    input [18:0] Wgt_9_385, // sfix19_En18 
    input [18:0] Wgt_9_386, // sfix19_En18 
    input [18:0] Wgt_9_387, // sfix19_En18 
    input [18:0] Wgt_9_388, // sfix19_En18 
    input [18:0] Wgt_9_389, // sfix19_En18 
    input [18:0] Wgt_9_390, // sfix19_En18 
    input [18:0] Wgt_9_391, // sfix19_En18 
    input [18:0] Wgt_9_392, // sfix19_En18 
    input [18:0] Wgt_9_393, // sfix19_En18 
    input [18:0] Wgt_9_394, // sfix19_En18 
    input [18:0] Wgt_9_395, // sfix19_En18 
    input [18:0] Wgt_9_396, // sfix19_En18 
    input [18:0] Wgt_9_397, // sfix19_En18 
    input [18:0] Wgt_9_398, // sfix19_En18 
    input [18:0] Wgt_9_399, // sfix19_En18 
    input [18:0] Wgt_9_400, // sfix19_En18 
    input [18:0] Wgt_9_401, // sfix19_En18 
    input [18:0] Wgt_9_402, // sfix19_En18 
    input [18:0] Wgt_9_403, // sfix19_En18 
    input [18:0] Wgt_9_404, // sfix19_En18 
    input [18:0] Wgt_9_405, // sfix19_En18 
    input [18:0] Wgt_9_406, // sfix19_En18 
    input [18:0] Wgt_9_407, // sfix19_En18 
    input [18:0] Wgt_9_408, // sfix19_En18 
    input [18:0] Wgt_9_409, // sfix19_En18 
    input [18:0] Wgt_9_410, // sfix19_En18 
    input [18:0] Wgt_9_411, // sfix19_En18 
    input [18:0] Wgt_9_412, // sfix19_En18 
    input [18:0] Wgt_9_413, // sfix19_En18 
    input [18:0] Wgt_9_414, // sfix19_En18 
    input [18:0] Wgt_9_415, // sfix19_En18 
    input [18:0] Wgt_9_416, // sfix19_En18 
    input [18:0] Wgt_9_417, // sfix19_En18 
    input [18:0] Wgt_9_418, // sfix19_En18 
    input [18:0] Wgt_9_419, // sfix19_En18 
    input [18:0] Wgt_9_420, // sfix19_En18 
    input [18:0] Wgt_9_421, // sfix19_En18 
    input [18:0] Wgt_9_422, // sfix19_En18 
    input [18:0] Wgt_9_423, // sfix19_En18 
    input [18:0] Wgt_9_424, // sfix19_En18 
    input [18:0] Wgt_9_425, // sfix19_En18 
    input [18:0] Wgt_9_426, // sfix19_En18 
    input [18:0] Wgt_9_427, // sfix19_En18 
    input [18:0] Wgt_9_428, // sfix19_En18 
    input [18:0] Wgt_9_429, // sfix19_En18 
    input [18:0] Wgt_9_430, // sfix19_En18 
    input [18:0] Wgt_9_431, // sfix19_En18 
    input [18:0] Wgt_9_432, // sfix19_En18 
    input [18:0] Wgt_9_433, // sfix19_En18 
    input [18:0] Wgt_9_434, // sfix19_En18 
    input [18:0] Wgt_9_435, // sfix19_En18 
    input [18:0] Wgt_9_436, // sfix19_En18 
    input [18:0] Wgt_9_437, // sfix19_En18 
    input [18:0] Wgt_9_438, // sfix19_En18 
    input [18:0] Wgt_9_439, // sfix19_En18 
    input [18:0] Wgt_9_440, // sfix19_En18 
    input [18:0] Wgt_9_441, // sfix19_En18 
    input [18:0] Wgt_9_442, // sfix19_En18 
    input [18:0] Wgt_9_443, // sfix19_En18 
    input [18:0] Wgt_9_444, // sfix19_En18 
    input [18:0] Wgt_9_445, // sfix19_En18 
    input [18:0] Wgt_9_446, // sfix19_En18 
    input [18:0] Wgt_9_447, // sfix19_En18 
    input [18:0] Wgt_9_448, // sfix19_En18 
    input [18:0] Wgt_9_449, // sfix19_En18 
    input [18:0] Wgt_9_450, // sfix19_En18 
    input [18:0] Wgt_9_451, // sfix19_En18 
    input [18:0] Wgt_9_452, // sfix19_En18 
    input [18:0] Wgt_9_453, // sfix19_En18 
    input [18:0] Wgt_9_454, // sfix19_En18 
    input [18:0] Wgt_9_455, // sfix19_En18 
    input [18:0] Wgt_9_456, // sfix19_En18 
    input [18:0] Wgt_9_457, // sfix19_En18 
    input [18:0] Wgt_9_458, // sfix19_En18 
    input [18:0] Wgt_9_459, // sfix19_En18 
    input [18:0] Wgt_9_460, // sfix19_En18 
    input [18:0] Wgt_9_461, // sfix19_En18 
    input [18:0] Wgt_9_462, // sfix19_En18 
    input [18:0] Wgt_9_463, // sfix19_En18 
    input [18:0] Wgt_9_464, // sfix19_En18 
    input [18:0] Wgt_9_465, // sfix19_En18 
    input [18:0] Wgt_9_466, // sfix19_En18 
    input [18:0] Wgt_9_467, // sfix19_En18 
    input [18:0] Wgt_9_468, // sfix19_En18 
    input [18:0] Wgt_9_469, // sfix19_En18 
    input [18:0] Wgt_9_470, // sfix19_En18 
    input [18:0] Wgt_9_471, // sfix19_En18 
    input [18:0] Wgt_9_472, // sfix19_En18 
    input [18:0] Wgt_9_473, // sfix19_En18 
    input [18:0] Wgt_9_474, // sfix19_En18 
    input [18:0] Wgt_9_475, // sfix19_En18 
    input [18:0] Wgt_9_476, // sfix19_En18 
    input [18:0] Wgt_9_477, // sfix19_En18 
    input [18:0] Wgt_9_478, // sfix19_En18 
    input [18:0] Wgt_9_479, // sfix19_En18 
    input [18:0] Wgt_9_480, // sfix19_En18 
    input [18:0] Wgt_9_481, // sfix19_En18 
    input [18:0] Wgt_9_482, // sfix19_En18 
    input [18:0] Wgt_9_483, // sfix19_En18 
    input [18:0] Wgt_9_484, // sfix19_En18 
    input [18:0] Wgt_9_485, // sfix19_En18 
    input [18:0] Wgt_9_486, // sfix19_En18 
    input [18:0] Wgt_9_487, // sfix19_En18 
    input [18:0] Wgt_9_488, // sfix19_En18 
    input [18:0] Wgt_9_489, // sfix19_En18 
    input [18:0] Wgt_9_490, // sfix19_En18 
    input [18:0] Wgt_9_491, // sfix19_En18 
    input [18:0] Wgt_9_492, // sfix19_En18 
    input [18:0] Wgt_9_493, // sfix19_En18 
    input [18:0] Wgt_9_494, // sfix19_En18 
    input [18:0] Wgt_9_495, // sfix19_En18 
    input [18:0] Wgt_9_496, // sfix19_En18 
    input [18:0] Wgt_9_497, // sfix19_En18 
    input [18:0] Wgt_9_498, // sfix19_En18 
    input [18:0] Wgt_9_499, // sfix19_En18 
    input [18:0] Wgt_9_500, // sfix19_En18 
    input [18:0] Wgt_9_501, // sfix19_En18 
    input [18:0] Wgt_9_502, // sfix19_En18 
    input [18:0] Wgt_9_503, // sfix19_En18 
    input [18:0] Wgt_9_504, // sfix19_En18 
    input [18:0] Wgt_9_505, // sfix19_En18 
    input [18:0] Wgt_9_506, // sfix19_En18 
    input [18:0] Wgt_9_507, // sfix19_En18 
    input [18:0] Wgt_9_508, // sfix19_En18 
    input [18:0] Wgt_9_509, // sfix19_En18 
    input [18:0] Wgt_9_510, // sfix19_En18 
    input [18:0] Wgt_9_511, // sfix19_En18 
    input [18:0] Wgt_9_512, // sfix19_En18 
    input [18:0] Wgt_9_513, // sfix19_En18 
    input [18:0] Wgt_9_514, // sfix19_En18 
    input [18:0] Wgt_9_515, // sfix19_En18 
    input [18:0] Wgt_9_516, // sfix19_En18 
    input [18:0] Wgt_9_517, // sfix19_En18 
    input [18:0] Wgt_9_518, // sfix19_En18 
    input [18:0] Wgt_9_519, // sfix19_En18 
    input [18:0] Wgt_9_520, // sfix19_En18 
    input [18:0] Wgt_9_521, // sfix19_En18 
    input [18:0] Wgt_9_522, // sfix19_En18 
    input [18:0] Wgt_9_523, // sfix19_En18 
    input [18:0] Wgt_9_524, // sfix19_En18 
    input [18:0] Wgt_9_525, // sfix19_En18 
    input [18:0] Wgt_9_526, // sfix19_En18 
    input [18:0] Wgt_9_527, // sfix19_En18 
    input [18:0] Wgt_9_528, // sfix19_En18 
    input [18:0] Wgt_9_529, // sfix19_En18 
    input [18:0] Wgt_9_530, // sfix19_En18 
    input [18:0] Wgt_9_531, // sfix19_En18 
    input [18:0] Wgt_9_532, // sfix19_En18 
    input [18:0] Wgt_9_533, // sfix19_En18 
    input [18:0] Wgt_9_534, // sfix19_En18 
    input [18:0] Wgt_9_535, // sfix19_En18 
    input [18:0] Wgt_9_536, // sfix19_En18 
    input [18:0] Wgt_9_537, // sfix19_En18 
    input [18:0] Wgt_9_538, // sfix19_En18 
    input [18:0] Wgt_9_539, // sfix19_En18 
    input [18:0] Wgt_9_540, // sfix19_En18 
    input [18:0] Wgt_9_541, // sfix19_En18 
    input [18:0] Wgt_9_542, // sfix19_En18 
    input [18:0] Wgt_9_543, // sfix19_En18 
    input [18:0] Wgt_9_544, // sfix19_En18 
    input [18:0] Wgt_9_545, // sfix19_En18 
    input [18:0] Wgt_9_546, // sfix19_En18 
    input [18:0] Wgt_9_547, // sfix19_En18 
    input [18:0] Wgt_9_548, // sfix19_En18 
    input [18:0] Wgt_9_549, // sfix19_En18 
    input [18:0] Wgt_9_550, // sfix19_En18 
    input [18:0] Wgt_9_551, // sfix19_En18 
    input [18:0] Wgt_9_552, // sfix19_En18 
    input [18:0] Wgt_9_553, // sfix19_En18 
    input [18:0] Wgt_9_554, // sfix19_En18 
    input [18:0] Wgt_9_555, // sfix19_En18 
    input [18:0] Wgt_9_556, // sfix19_En18 
    input [18:0] Wgt_9_557, // sfix19_En18 
    input [18:0] Wgt_9_558, // sfix19_En18 
    input [18:0] Wgt_9_559, // sfix19_En18 
    input [18:0] Wgt_9_560, // sfix19_En18 
    input [18:0] Wgt_9_561, // sfix19_En18 
    input [18:0] Wgt_9_562, // sfix19_En18 
    input [18:0] Wgt_9_563, // sfix19_En18 
    input [18:0] Wgt_9_564, // sfix19_En18 
    input [18:0] Wgt_9_565, // sfix19_En18 
    input [18:0] Wgt_9_566, // sfix19_En18 
    input [18:0] Wgt_9_567, // sfix19_En18 
    input [18:0] Wgt_9_568, // sfix19_En18 
    input [18:0] Wgt_9_569, // sfix19_En18 
    input [18:0] Wgt_9_570, // sfix19_En18 
    input [18:0] Wgt_9_571, // sfix19_En18 
    input [18:0] Wgt_9_572, // sfix19_En18 
    input [18:0] Wgt_9_573, // sfix19_En18 
    input [18:0] Wgt_9_574, // sfix19_En18 
    input [18:0] Wgt_9_575, // sfix19_En18 
    input [18:0] Wgt_9_576, // sfix19_En18 
    input [18:0] Wgt_9_577, // sfix19_En18 
    input [18:0] Wgt_9_578, // sfix19_En18 
    input [18:0] Wgt_9_579, // sfix19_En18 
    input [18:0] Wgt_9_580, // sfix19_En18 
    input [18:0] Wgt_9_581, // sfix19_En18 
    input [18:0] Wgt_9_582, // sfix19_En18 
    input [18:0] Wgt_9_583, // sfix19_En18 
    input [18:0] Wgt_9_584, // sfix19_En18 
    input [18:0] Wgt_9_585, // sfix19_En18 
    input [18:0] Wgt_9_586, // sfix19_En18 
    input [18:0] Wgt_9_587, // sfix19_En18 
    input [18:0] Wgt_9_588, // sfix19_En18 
    input [18:0] Wgt_9_589, // sfix19_En18 
    input [18:0] Wgt_9_590, // sfix19_En18 
    input [18:0] Wgt_9_591, // sfix19_En18 
    input [18:0] Wgt_9_592, // sfix19_En18 
    input [18:0] Wgt_9_593, // sfix19_En18 
    input [18:0] Wgt_9_594, // sfix19_En18 
    input [18:0] Wgt_9_595, // sfix19_En18 
    input [18:0] Wgt_9_596, // sfix19_En18 
    input [18:0] Wgt_9_597, // sfix19_En18 
    input [18:0] Wgt_9_598, // sfix19_En18 
    input [18:0] Wgt_9_599, // sfix19_En18 
    input [18:0] Wgt_9_600, // sfix19_En18 
    input [18:0] Wgt_9_601, // sfix19_En18 
    input [18:0] Wgt_9_602, // sfix19_En18 
    input [18:0] Wgt_9_603, // sfix19_En18 
    input [18:0] Wgt_9_604, // sfix19_En18 
    input [18:0] Wgt_9_605, // sfix19_En18 
    input [18:0] Wgt_9_606, // sfix19_En18 
    input [18:0] Wgt_9_607, // sfix19_En18 
    input [18:0] Wgt_9_608, // sfix19_En18 
    input [18:0] Wgt_9_609, // sfix19_En18 
    input [18:0] Wgt_9_610, // sfix19_En18 
    input [18:0] Wgt_9_611, // sfix19_En18 
    input [18:0] Wgt_9_612, // sfix19_En18 
    input [18:0] Wgt_9_613, // sfix19_En18 
    input [18:0] Wgt_9_614, // sfix19_En18 
    input [18:0] Wgt_9_615, // sfix19_En18 
    input [18:0] Wgt_9_616, // sfix19_En18 
    input [18:0] Wgt_9_617, // sfix19_En18 
    input [18:0] Wgt_9_618, // sfix19_En18 
    input [18:0] Wgt_9_619, // sfix19_En18 
    input [18:0] Wgt_9_620, // sfix19_En18 
    input [18:0] Wgt_9_621, // sfix19_En18 
    input [18:0] Wgt_9_622, // sfix19_En18 
    input [18:0] Wgt_9_623, // sfix19_En18 
    input [18:0] Wgt_9_624, // sfix19_En18 
    input [18:0] Wgt_9_625, // sfix19_En18 
    input [18:0] Wgt_9_626, // sfix19_En18 
    input [18:0] Wgt_9_627, // sfix19_En18 
    input [18:0] Wgt_9_628, // sfix19_En18 
    input [18:0] Wgt_9_629, // sfix19_En18 
    input [18:0] Wgt_9_630, // sfix19_En18 
    input [18:0] Wgt_9_631, // sfix19_En18 
    input [18:0] Wgt_9_632, // sfix19_En18 
    input [18:0] Wgt_9_633, // sfix19_En18 
    input [18:0] Wgt_9_634, // sfix19_En18 
    input [18:0] Wgt_9_635, // sfix19_En18 
    input [18:0] Wgt_9_636, // sfix19_En18 
    input [18:0] Wgt_9_637, // sfix19_En18 
    input [18:0] Wgt_9_638, // sfix19_En18 
    input [18:0] Wgt_9_639, // sfix19_En18 
    input [18:0] Wgt_9_640, // sfix19_En18 
    input [18:0] Wgt_9_641, // sfix19_En18 
    input [18:0] Wgt_9_642, // sfix19_En18 
    input [18:0] Wgt_9_643, // sfix19_En18 
    input [18:0] Wgt_9_644, // sfix19_En18 
    input [18:0] Wgt_9_645, // sfix19_En18 
    input [18:0] Wgt_9_646, // sfix19_En18 
    input [18:0] Wgt_9_647, // sfix19_En18 
    input [18:0] Wgt_9_648, // sfix19_En18 
    input [18:0] Wgt_9_649, // sfix19_En18 
    input [18:0] Wgt_9_650, // sfix19_En18 
    input [18:0] Wgt_9_651, // sfix19_En18 
    input [18:0] Wgt_9_652, // sfix19_En18 
    input [18:0] Wgt_9_653, // sfix19_En18 
    input [18:0] Wgt_9_654, // sfix19_En18 
    input [18:0] Wgt_9_655, // sfix19_En18 
    input [18:0] Wgt_9_656, // sfix19_En18 
    input [18:0] Wgt_9_657, // sfix19_En18 
    input [18:0] Wgt_9_658, // sfix19_En18 
    input [18:0] Wgt_9_659, // sfix19_En18 
    input [18:0] Wgt_9_660, // sfix19_En18 
    input [18:0] Wgt_9_661, // sfix19_En18 
    input [18:0] Wgt_9_662, // sfix19_En18 
    input [18:0] Wgt_9_663, // sfix19_En18 
    input [18:0] Wgt_9_664, // sfix19_En18 
    input [18:0] Wgt_9_665, // sfix19_En18 
    input [18:0] Wgt_9_666, // sfix19_En18 
    input [18:0] Wgt_9_667, // sfix19_En18 
    input [18:0] Wgt_9_668, // sfix19_En18 
    input [18:0] Wgt_9_669, // sfix19_En18 
    input [18:0] Wgt_9_670, // sfix19_En18 
    input [18:0] Wgt_9_671, // sfix19_En18 
    input [18:0] Wgt_9_672, // sfix19_En18 
    input [18:0] Wgt_9_673, // sfix19_En18 
    input [18:0] Wgt_9_674, // sfix19_En18 
    input [18:0] Wgt_9_675, // sfix19_En18 
    input [18:0] Wgt_9_676, // sfix19_En18 
    input [18:0] Wgt_9_677, // sfix19_En18 
    input [18:0] Wgt_9_678, // sfix19_En18 
    input [18:0] Wgt_9_679, // sfix19_En18 
    input [18:0] Wgt_9_680, // sfix19_En18 
    input [18:0] Wgt_9_681, // sfix19_En18 
    input [18:0] Wgt_9_682, // sfix19_En18 
    input [18:0] Wgt_9_683, // sfix19_En18 
    input [18:0] Wgt_9_684, // sfix19_En18 
    input [18:0] Wgt_9_685, // sfix19_En18 
    input [18:0] Wgt_9_686, // sfix19_En18 
    input [18:0] Wgt_9_687, // sfix19_En18 
    input [18:0] Wgt_9_688, // sfix19_En18 
    input [18:0] Wgt_9_689, // sfix19_En18 
    input [18:0] Wgt_9_690, // sfix19_En18 
    input [18:0] Wgt_9_691, // sfix19_En18 
    input [18:0] Wgt_9_692, // sfix19_En18 
    input [18:0] Wgt_9_693, // sfix19_En18 
    input [18:0] Wgt_9_694, // sfix19_En18 
    input [18:0] Wgt_9_695, // sfix19_En18 
    input [18:0] Wgt_9_696, // sfix19_En18 
    input [18:0] Wgt_9_697, // sfix19_En18 
    input [18:0] Wgt_9_698, // sfix19_En18 
    input [18:0] Wgt_9_699, // sfix19_En18 
    input [18:0] Wgt_9_700, // sfix19_En18 
    input [18:0] Wgt_9_701, // sfix19_En18 
    input [18:0] Wgt_9_702, // sfix19_En18 
    input [18:0] Wgt_9_703, // sfix19_En18 
    input [18:0] Wgt_9_704, // sfix19_En18 
    input [18:0] Wgt_9_705, // sfix19_En18 
    input [18:0] Wgt_9_706, // sfix19_En18 
    input [18:0] Wgt_9_707, // sfix19_En18 
    input [18:0] Wgt_9_708, // sfix19_En18 
    input [18:0] Wgt_9_709, // sfix19_En18 
    input [18:0] Wgt_9_710, // sfix19_En18 
    input [18:0] Wgt_9_711, // sfix19_En18 
    input [18:0] Wgt_9_712, // sfix19_En18 
    input [18:0] Wgt_9_713, // sfix19_En18 
    input [18:0] Wgt_9_714, // sfix19_En18 
    input [18:0] Wgt_9_715, // sfix19_En18 
    input [18:0] Wgt_9_716, // sfix19_En18 
    input [18:0] Wgt_9_717, // sfix19_En18 
    input [18:0] Wgt_9_718, // sfix19_En18 
    input [18:0] Wgt_9_719, // sfix19_En18 
    input [18:0] Wgt_9_720, // sfix19_En18 
    input [18:0] Wgt_9_721, // sfix19_En18 
    input [18:0] Wgt_9_722, // sfix19_En18 
    input [18:0] Wgt_9_723, // sfix19_En18 
    input [18:0] Wgt_9_724, // sfix19_En18 
    input [18:0] Wgt_9_725, // sfix19_En18 
    input [18:0] Wgt_9_726, // sfix19_En18 
    input [18:0] Wgt_9_727, // sfix19_En18 
    input [18:0] Wgt_9_728, // sfix19_En18 
    input [18:0] Wgt_9_729, // sfix19_En18 
    input [18:0] Wgt_9_730, // sfix19_En18 
    input [18:0] Wgt_9_731, // sfix19_En18 
    input [18:0] Wgt_9_732, // sfix19_En18 
    input [18:0] Wgt_9_733, // sfix19_En18 
    input [18:0] Wgt_9_734, // sfix19_En18 
    input [18:0] Wgt_9_735, // sfix19_En18 
    input [18:0] Wgt_9_736, // sfix19_En18 
    input [18:0] Wgt_9_737, // sfix19_En18 
    input [18:0] Wgt_9_738, // sfix19_En18 
    input [18:0] Wgt_9_739, // sfix19_En18 
    input [18:0] Wgt_9_740, // sfix19_En18 
    input [18:0] Wgt_9_741, // sfix19_En18 
    input [18:0] Wgt_9_742, // sfix19_En18 
    input [18:0] Wgt_9_743, // sfix19_En18 
    input [18:0] Wgt_9_744, // sfix19_En18 
    input [18:0] Wgt_9_745, // sfix19_En18 
    input [18:0] Wgt_9_746, // sfix19_En18 
    input [18:0] Wgt_9_747, // sfix19_En18 
    input [18:0] Wgt_9_748, // sfix19_En18 
    input [18:0] Wgt_9_749, // sfix19_En18 
    input [18:0] Wgt_9_750, // sfix19_En18 
    input [18:0] Wgt_9_751, // sfix19_En18 
    input [18:0] Wgt_9_752, // sfix19_En18 
    input [18:0] Wgt_9_753, // sfix19_En18 
    input [18:0] Wgt_9_754, // sfix19_En18 
    input [18:0] Wgt_9_755, // sfix19_En18 
    input [18:0] Wgt_9_756, // sfix19_En18 
    input [18:0] Wgt_9_757, // sfix19_En18 
    input [18:0] Wgt_9_758, // sfix19_En18 
    input [18:0] Wgt_9_759, // sfix19_En18 
    input [18:0] Wgt_9_760, // sfix19_En18 
    input [18:0] Wgt_9_761, // sfix19_En18 
    input [18:0] Wgt_9_762, // sfix19_En18 
    input [18:0] Wgt_9_763, // sfix19_En18 
    input [18:0] Wgt_9_764, // sfix19_En18 
    input [18:0] Wgt_9_765, // sfix19_En18 
    input [18:0] Wgt_9_766, // sfix19_En18 
    input [18:0] Wgt_9_767, // sfix19_En18 
    input [18:0] Wgt_9_768, // sfix19_En18 
    input [18:0] Wgt_9_769, // sfix19_En18 
    input [18:0] Wgt_9_770, // sfix19_En18 
    input [18:0] Wgt_9_771, // sfix19_En18 
    input [18:0] Wgt_9_772, // sfix19_En18 
    input [18:0] Wgt_9_773, // sfix19_En18 
    input [18:0] Wgt_9_774, // sfix19_En18 
    input [18:0] Wgt_9_775, // sfix19_En18 
    input [18:0] Wgt_9_776, // sfix19_En18 
    input [18:0] Wgt_9_777, // sfix19_En18 
    input [18:0] Wgt_9_778, // sfix19_En18 
    input [18:0] Wgt_9_779, // sfix19_En18 
    input [18:0] Wgt_9_780, // sfix19_En18 
    input [18:0] Wgt_9_781, // sfix19_En18 
    input [18:0] Wgt_9_782, // sfix19_En18 
    input [18:0] Wgt_9_783, // sfix19_En18 
    input [18:0] Wgt_9_784, // sfix19_En18 
    input [9:0] Pix_0, // sfix10_En0 
    input [9:0] Pix_1, // sfix10_En0 
    input [9:0] Pix_2, // sfix10_En0 
    input [9:0] Pix_3, // sfix10_En0 
    input [9:0] Pix_4, // sfix10_En0 
    input [9:0] Pix_5, // sfix10_En0 
    input [9:0] Pix_6, // sfix10_En0 
    input [9:0] Pix_7, // sfix10_En0 
    input [9:0] Pix_8, // sfix10_En0 
    input [9:0] Pix_9, // sfix10_En0 
    input [9:0] Pix_10, // sfix10_En0 
    input [9:0] Pix_11, // sfix10_En0 
    input [9:0] Pix_12, // sfix10_En0 
    input [9:0] Pix_13, // sfix10_En0 
    input [9:0] Pix_14, // sfix10_En0 
    input [9:0] Pix_15, // sfix10_En0 
    input [9:0] Pix_16, // sfix10_En0 
    input [9:0] Pix_17, // sfix10_En0 
    input [9:0] Pix_18, // sfix10_En0 
    input [9:0] Pix_19, // sfix10_En0 
    input [9:0] Pix_20, // sfix10_En0 
    input [9:0] Pix_21, // sfix10_En0 
    input [9:0] Pix_22, // sfix10_En0 
    input [9:0] Pix_23, // sfix10_En0 
    input [9:0] Pix_24, // sfix10_En0 
    input [9:0] Pix_25, // sfix10_En0 
    input [9:0] Pix_26, // sfix10_En0 
    input [9:0] Pix_27, // sfix10_En0 
    input [9:0] Pix_28, // sfix10_En0 
    input [9:0] Pix_29, // sfix10_En0 
    input [9:0] Pix_30, // sfix10_En0 
    input [9:0] Pix_31, // sfix10_En0 
    input [9:0] Pix_32, // sfix10_En0 
    input [9:0] Pix_33, // sfix10_En0 
    input [9:0] Pix_34, // sfix10_En0 
    input [9:0] Pix_35, // sfix10_En0 
    input [9:0] Pix_36, // sfix10_En0 
    input [9:0] Pix_37, // sfix10_En0 
    input [9:0] Pix_38, // sfix10_En0 
    input [9:0] Pix_39, // sfix10_En0 
    input [9:0] Pix_40, // sfix10_En0 
    input [9:0] Pix_41, // sfix10_En0 
    input [9:0] Pix_42, // sfix10_En0 
    input [9:0] Pix_43, // sfix10_En0 
    input [9:0] Pix_44, // sfix10_En0 
    input [9:0] Pix_45, // sfix10_En0 
    input [9:0] Pix_46, // sfix10_En0 
    input [9:0] Pix_47, // sfix10_En0 
    input [9:0] Pix_48, // sfix10_En0 
    input [9:0] Pix_49, // sfix10_En0 
    input [9:0] Pix_50, // sfix10_En0 
    input [9:0] Pix_51, // sfix10_En0 
    input [9:0] Pix_52, // sfix10_En0 
    input [9:0] Pix_53, // sfix10_En0 
    input [9:0] Pix_54, // sfix10_En0 
    input [9:0] Pix_55, // sfix10_En0 
    input [9:0] Pix_56, // sfix10_En0 
    input [9:0] Pix_57, // sfix10_En0 
    input [9:0] Pix_58, // sfix10_En0 
    input [9:0] Pix_59, // sfix10_En0 
    input [9:0] Pix_60, // sfix10_En0 
    input [9:0] Pix_61, // sfix10_En0 
    input [9:0] Pix_62, // sfix10_En0 
    input [9:0] Pix_63, // sfix10_En0 
    input [9:0] Pix_64, // sfix10_En0 
    input [9:0] Pix_65, // sfix10_En0 
    input [9:0] Pix_66, // sfix10_En0 
    input [9:0] Pix_67, // sfix10_En0 
    input [9:0] Pix_68, // sfix10_En0 
    input [9:0] Pix_69, // sfix10_En0 
    input [9:0] Pix_70, // sfix10_En0 
    input [9:0] Pix_71, // sfix10_En0 
    input [9:0] Pix_72, // sfix10_En0 
    input [9:0] Pix_73, // sfix10_En0 
    input [9:0] Pix_74, // sfix10_En0 
    input [9:0] Pix_75, // sfix10_En0 
    input [9:0] Pix_76, // sfix10_En0 
    input [9:0] Pix_77, // sfix10_En0 
    input [9:0] Pix_78, // sfix10_En0 
    input [9:0] Pix_79, // sfix10_En0 
    input [9:0] Pix_80, // sfix10_En0 
    input [9:0] Pix_81, // sfix10_En0 
    input [9:0] Pix_82, // sfix10_En0 
    input [9:0] Pix_83, // sfix10_En0 
    input [9:0] Pix_84, // sfix10_En0 
    input [9:0] Pix_85, // sfix10_En0 
    input [9:0] Pix_86, // sfix10_En0 
    input [9:0] Pix_87, // sfix10_En0 
    input [9:0] Pix_88, // sfix10_En0 
    input [9:0] Pix_89, // sfix10_En0 
    input [9:0] Pix_90, // sfix10_En0 
    input [9:0] Pix_91, // sfix10_En0 
    input [9:0] Pix_92, // sfix10_En0 
    input [9:0] Pix_93, // sfix10_En0 
    input [9:0] Pix_94, // sfix10_En0 
    input [9:0] Pix_95, // sfix10_En0 
    input [9:0] Pix_96, // sfix10_En0 
    input [9:0] Pix_97, // sfix10_En0 
    input [9:0] Pix_98, // sfix10_En0 
    input [9:0] Pix_99, // sfix10_En0 
    input [9:0] Pix_100, // sfix10_En0 
    input [9:0] Pix_101, // sfix10_En0 
    input [9:0] Pix_102, // sfix10_En0 
    input [9:0] Pix_103, // sfix10_En0 
    input [9:0] Pix_104, // sfix10_En0 
    input [9:0] Pix_105, // sfix10_En0 
    input [9:0] Pix_106, // sfix10_En0 
    input [9:0] Pix_107, // sfix10_En0 
    input [9:0] Pix_108, // sfix10_En0 
    input [9:0] Pix_109, // sfix10_En0 
    input [9:0] Pix_110, // sfix10_En0 
    input [9:0] Pix_111, // sfix10_En0 
    input [9:0] Pix_112, // sfix10_En0 
    input [9:0] Pix_113, // sfix10_En0 
    input [9:0] Pix_114, // sfix10_En0 
    input [9:0] Pix_115, // sfix10_En0 
    input [9:0] Pix_116, // sfix10_En0 
    input [9:0] Pix_117, // sfix10_En0 
    input [9:0] Pix_118, // sfix10_En0 
    input [9:0] Pix_119, // sfix10_En0 
    input [9:0] Pix_120, // sfix10_En0 
    input [9:0] Pix_121, // sfix10_En0 
    input [9:0] Pix_122, // sfix10_En0 
    input [9:0] Pix_123, // sfix10_En0 
    input [9:0] Pix_124, // sfix10_En0 
    input [9:0] Pix_125, // sfix10_En0 
    input [9:0] Pix_126, // sfix10_En0 
    input [9:0] Pix_127, // sfix10_En0 
    input [9:0] Pix_128, // sfix10_En0 
    input [9:0] Pix_129, // sfix10_En0 
    input [9:0] Pix_130, // sfix10_En0 
    input [9:0] Pix_131, // sfix10_En0 
    input [9:0] Pix_132, // sfix10_En0 
    input [9:0] Pix_133, // sfix10_En0 
    input [9:0] Pix_134, // sfix10_En0 
    input [9:0] Pix_135, // sfix10_En0 
    input [9:0] Pix_136, // sfix10_En0 
    input [9:0] Pix_137, // sfix10_En0 
    input [9:0] Pix_138, // sfix10_En0 
    input [9:0] Pix_139, // sfix10_En0 
    input [9:0] Pix_140, // sfix10_En0 
    input [9:0] Pix_141, // sfix10_En0 
    input [9:0] Pix_142, // sfix10_En0 
    input [9:0] Pix_143, // sfix10_En0 
    input [9:0] Pix_144, // sfix10_En0 
    input [9:0] Pix_145, // sfix10_En0 
    input [9:0] Pix_146, // sfix10_En0 
    input [9:0] Pix_147, // sfix10_En0 
    input [9:0] Pix_148, // sfix10_En0 
    input [9:0] Pix_149, // sfix10_En0 
    input [9:0] Pix_150, // sfix10_En0 
    input [9:0] Pix_151, // sfix10_En0 
    input [9:0] Pix_152, // sfix10_En0 
    input [9:0] Pix_153, // sfix10_En0 
    input [9:0] Pix_154, // sfix10_En0 
    input [9:0] Pix_155, // sfix10_En0 
    input [9:0] Pix_156, // sfix10_En0 
    input [9:0] Pix_157, // sfix10_En0 
    input [9:0] Pix_158, // sfix10_En0 
    input [9:0] Pix_159, // sfix10_En0 
    input [9:0] Pix_160, // sfix10_En0 
    input [9:0] Pix_161, // sfix10_En0 
    input [9:0] Pix_162, // sfix10_En0 
    input [9:0] Pix_163, // sfix10_En0 
    input [9:0] Pix_164, // sfix10_En0 
    input [9:0] Pix_165, // sfix10_En0 
    input [9:0] Pix_166, // sfix10_En0 
    input [9:0] Pix_167, // sfix10_En0 
    input [9:0] Pix_168, // sfix10_En0 
    input [9:0] Pix_169, // sfix10_En0 
    input [9:0] Pix_170, // sfix10_En0 
    input [9:0] Pix_171, // sfix10_En0 
    input [9:0] Pix_172, // sfix10_En0 
    input [9:0] Pix_173, // sfix10_En0 
    input [9:0] Pix_174, // sfix10_En0 
    input [9:0] Pix_175, // sfix10_En0 
    input [9:0] Pix_176, // sfix10_En0 
    input [9:0] Pix_177, // sfix10_En0 
    input [9:0] Pix_178, // sfix10_En0 
    input [9:0] Pix_179, // sfix10_En0 
    input [9:0] Pix_180, // sfix10_En0 
    input [9:0] Pix_181, // sfix10_En0 
    input [9:0] Pix_182, // sfix10_En0 
    input [9:0] Pix_183, // sfix10_En0 
    input [9:0] Pix_184, // sfix10_En0 
    input [9:0] Pix_185, // sfix10_En0 
    input [9:0] Pix_186, // sfix10_En0 
    input [9:0] Pix_187, // sfix10_En0 
    input [9:0] Pix_188, // sfix10_En0 
    input [9:0] Pix_189, // sfix10_En0 
    input [9:0] Pix_190, // sfix10_En0 
    input [9:0] Pix_191, // sfix10_En0 
    input [9:0] Pix_192, // sfix10_En0 
    input [9:0] Pix_193, // sfix10_En0 
    input [9:0] Pix_194, // sfix10_En0 
    input [9:0] Pix_195, // sfix10_En0 
    input [9:0] Pix_196, // sfix10_En0 
    input [9:0] Pix_197, // sfix10_En0 
    input [9:0] Pix_198, // sfix10_En0 
    input [9:0] Pix_199, // sfix10_En0 
    input [9:0] Pix_200, // sfix10_En0 
    input [9:0] Pix_201, // sfix10_En0 
    input [9:0] Pix_202, // sfix10_En0 
    input [9:0] Pix_203, // sfix10_En0 
    input [9:0] Pix_204, // sfix10_En0 
    input [9:0] Pix_205, // sfix10_En0 
    input [9:0] Pix_206, // sfix10_En0 
    input [9:0] Pix_207, // sfix10_En0 
    input [9:0] Pix_208, // sfix10_En0 
    input [9:0] Pix_209, // sfix10_En0 
    input [9:0] Pix_210, // sfix10_En0 
    input [9:0] Pix_211, // sfix10_En0 
    input [9:0] Pix_212, // sfix10_En0 
    input [9:0] Pix_213, // sfix10_En0 
    input [9:0] Pix_214, // sfix10_En0 
    input [9:0] Pix_215, // sfix10_En0 
    input [9:0] Pix_216, // sfix10_En0 
    input [9:0] Pix_217, // sfix10_En0 
    input [9:0] Pix_218, // sfix10_En0 
    input [9:0] Pix_219, // sfix10_En0 
    input [9:0] Pix_220, // sfix10_En0 
    input [9:0] Pix_221, // sfix10_En0 
    input [9:0] Pix_222, // sfix10_En0 
    input [9:0] Pix_223, // sfix10_En0 
    input [9:0] Pix_224, // sfix10_En0 
    input [9:0] Pix_225, // sfix10_En0 
    input [9:0] Pix_226, // sfix10_En0 
    input [9:0] Pix_227, // sfix10_En0 
    input [9:0] Pix_228, // sfix10_En0 
    input [9:0] Pix_229, // sfix10_En0 
    input [9:0] Pix_230, // sfix10_En0 
    input [9:0] Pix_231, // sfix10_En0 
    input [9:0] Pix_232, // sfix10_En0 
    input [9:0] Pix_233, // sfix10_En0 
    input [9:0] Pix_234, // sfix10_En0 
    input [9:0] Pix_235, // sfix10_En0 
    input [9:0] Pix_236, // sfix10_En0 
    input [9:0] Pix_237, // sfix10_En0 
    input [9:0] Pix_238, // sfix10_En0 
    input [9:0] Pix_239, // sfix10_En0 
    input [9:0] Pix_240, // sfix10_En0 
    input [9:0] Pix_241, // sfix10_En0 
    input [9:0] Pix_242, // sfix10_En0 
    input [9:0] Pix_243, // sfix10_En0 
    input [9:0] Pix_244, // sfix10_En0 
    input [9:0] Pix_245, // sfix10_En0 
    input [9:0] Pix_246, // sfix10_En0 
    input [9:0] Pix_247, // sfix10_En0 
    input [9:0] Pix_248, // sfix10_En0 
    input [9:0] Pix_249, // sfix10_En0 
    input [9:0] Pix_250, // sfix10_En0 
    input [9:0] Pix_251, // sfix10_En0 
    input [9:0] Pix_252, // sfix10_En0 
    input [9:0] Pix_253, // sfix10_En0 
    input [9:0] Pix_254, // sfix10_En0 
    input [9:0] Pix_255, // sfix10_En0 
    input [9:0] Pix_256, // sfix10_En0 
    input [9:0] Pix_257, // sfix10_En0 
    input [9:0] Pix_258, // sfix10_En0 
    input [9:0] Pix_259, // sfix10_En0 
    input [9:0] Pix_260, // sfix10_En0 
    input [9:0] Pix_261, // sfix10_En0 
    input [9:0] Pix_262, // sfix10_En0 
    input [9:0] Pix_263, // sfix10_En0 
    input [9:0] Pix_264, // sfix10_En0 
    input [9:0] Pix_265, // sfix10_En0 
    input [9:0] Pix_266, // sfix10_En0 
    input [9:0] Pix_267, // sfix10_En0 
    input [9:0] Pix_268, // sfix10_En0 
    input [9:0] Pix_269, // sfix10_En0 
    input [9:0] Pix_270, // sfix10_En0 
    input [9:0] Pix_271, // sfix10_En0 
    input [9:0] Pix_272, // sfix10_En0 
    input [9:0] Pix_273, // sfix10_En0 
    input [9:0] Pix_274, // sfix10_En0 
    input [9:0] Pix_275, // sfix10_En0 
    input [9:0] Pix_276, // sfix10_En0 
    input [9:0] Pix_277, // sfix10_En0 
    input [9:0] Pix_278, // sfix10_En0 
    input [9:0] Pix_279, // sfix10_En0 
    input [9:0] Pix_280, // sfix10_En0 
    input [9:0] Pix_281, // sfix10_En0 
    input [9:0] Pix_282, // sfix10_En0 
    input [9:0] Pix_283, // sfix10_En0 
    input [9:0] Pix_284, // sfix10_En0 
    input [9:0] Pix_285, // sfix10_En0 
    input [9:0] Pix_286, // sfix10_En0 
    input [9:0] Pix_287, // sfix10_En0 
    input [9:0] Pix_288, // sfix10_En0 
    input [9:0] Pix_289, // sfix10_En0 
    input [9:0] Pix_290, // sfix10_En0 
    input [9:0] Pix_291, // sfix10_En0 
    input [9:0] Pix_292, // sfix10_En0 
    input [9:0] Pix_293, // sfix10_En0 
    input [9:0] Pix_294, // sfix10_En0 
    input [9:0] Pix_295, // sfix10_En0 
    input [9:0] Pix_296, // sfix10_En0 
    input [9:0] Pix_297, // sfix10_En0 
    input [9:0] Pix_298, // sfix10_En0 
    input [9:0] Pix_299, // sfix10_En0 
    input [9:0] Pix_300, // sfix10_En0 
    input [9:0] Pix_301, // sfix10_En0 
    input [9:0] Pix_302, // sfix10_En0 
    input [9:0] Pix_303, // sfix10_En0 
    input [9:0] Pix_304, // sfix10_En0 
    input [9:0] Pix_305, // sfix10_En0 
    input [9:0] Pix_306, // sfix10_En0 
    input [9:0] Pix_307, // sfix10_En0 
    input [9:0] Pix_308, // sfix10_En0 
    input [9:0] Pix_309, // sfix10_En0 
    input [9:0] Pix_310, // sfix10_En0 
    input [9:0] Pix_311, // sfix10_En0 
    input [9:0] Pix_312, // sfix10_En0 
    input [9:0] Pix_313, // sfix10_En0 
    input [9:0] Pix_314, // sfix10_En0 
    input [9:0] Pix_315, // sfix10_En0 
    input [9:0] Pix_316, // sfix10_En0 
    input [9:0] Pix_317, // sfix10_En0 
    input [9:0] Pix_318, // sfix10_En0 
    input [9:0] Pix_319, // sfix10_En0 
    input [9:0] Pix_320, // sfix10_En0 
    input [9:0] Pix_321, // sfix10_En0 
    input [9:0] Pix_322, // sfix10_En0 
    input [9:0] Pix_323, // sfix10_En0 
    input [9:0] Pix_324, // sfix10_En0 
    input [9:0] Pix_325, // sfix10_En0 
    input [9:0] Pix_326, // sfix10_En0 
    input [9:0] Pix_327, // sfix10_En0 
    input [9:0] Pix_328, // sfix10_En0 
    input [9:0] Pix_329, // sfix10_En0 
    input [9:0] Pix_330, // sfix10_En0 
    input [9:0] Pix_331, // sfix10_En0 
    input [9:0] Pix_332, // sfix10_En0 
    input [9:0] Pix_333, // sfix10_En0 
    input [9:0] Pix_334, // sfix10_En0 
    input [9:0] Pix_335, // sfix10_En0 
    input [9:0] Pix_336, // sfix10_En0 
    input [9:0] Pix_337, // sfix10_En0 
    input [9:0] Pix_338, // sfix10_En0 
    input [9:0] Pix_339, // sfix10_En0 
    input [9:0] Pix_340, // sfix10_En0 
    input [9:0] Pix_341, // sfix10_En0 
    input [9:0] Pix_342, // sfix10_En0 
    input [9:0] Pix_343, // sfix10_En0 
    input [9:0] Pix_344, // sfix10_En0 
    input [9:0] Pix_345, // sfix10_En0 
    input [9:0] Pix_346, // sfix10_En0 
    input [9:0] Pix_347, // sfix10_En0 
    input [9:0] Pix_348, // sfix10_En0 
    input [9:0] Pix_349, // sfix10_En0 
    input [9:0] Pix_350, // sfix10_En0 
    input [9:0] Pix_351, // sfix10_En0 
    input [9:0] Pix_352, // sfix10_En0 
    input [9:0] Pix_353, // sfix10_En0 
    input [9:0] Pix_354, // sfix10_En0 
    input [9:0] Pix_355, // sfix10_En0 
    input [9:0] Pix_356, // sfix10_En0 
    input [9:0] Pix_357, // sfix10_En0 
    input [9:0] Pix_358, // sfix10_En0 
    input [9:0] Pix_359, // sfix10_En0 
    input [9:0] Pix_360, // sfix10_En0 
    input [9:0] Pix_361, // sfix10_En0 
    input [9:0] Pix_362, // sfix10_En0 
    input [9:0] Pix_363, // sfix10_En0 
    input [9:0] Pix_364, // sfix10_En0 
    input [9:0] Pix_365, // sfix10_En0 
    input [9:0] Pix_366, // sfix10_En0 
    input [9:0] Pix_367, // sfix10_En0 
    input [9:0] Pix_368, // sfix10_En0 
    input [9:0] Pix_369, // sfix10_En0 
    input [9:0] Pix_370, // sfix10_En0 
    input [9:0] Pix_371, // sfix10_En0 
    input [9:0] Pix_372, // sfix10_En0 
    input [9:0] Pix_373, // sfix10_En0 
    input [9:0] Pix_374, // sfix10_En0 
    input [9:0] Pix_375, // sfix10_En0 
    input [9:0] Pix_376, // sfix10_En0 
    input [9:0] Pix_377, // sfix10_En0 
    input [9:0] Pix_378, // sfix10_En0 
    input [9:0] Pix_379, // sfix10_En0 
    input [9:0] Pix_380, // sfix10_En0 
    input [9:0] Pix_381, // sfix10_En0 
    input [9:0] Pix_382, // sfix10_En0 
    input [9:0] Pix_383, // sfix10_En0 
    input [9:0] Pix_384, // sfix10_En0 
    input [9:0] Pix_385, // sfix10_En0 
    input [9:0] Pix_386, // sfix10_En0 
    input [9:0] Pix_387, // sfix10_En0 
    input [9:0] Pix_388, // sfix10_En0 
    input [9:0] Pix_389, // sfix10_En0 
    input [9:0] Pix_390, // sfix10_En0 
    input [9:0] Pix_391, // sfix10_En0 
    input [9:0] Pix_392, // sfix10_En0 
    input [9:0] Pix_393, // sfix10_En0 
    input [9:0] Pix_394, // sfix10_En0 
    input [9:0] Pix_395, // sfix10_En0 
    input [9:0] Pix_396, // sfix10_En0 
    input [9:0] Pix_397, // sfix10_En0 
    input [9:0] Pix_398, // sfix10_En0 
    input [9:0] Pix_399, // sfix10_En0 
    input [9:0] Pix_400, // sfix10_En0 
    input [9:0] Pix_401, // sfix10_En0 
    input [9:0] Pix_402, // sfix10_En0 
    input [9:0] Pix_403, // sfix10_En0 
    input [9:0] Pix_404, // sfix10_En0 
    input [9:0] Pix_405, // sfix10_En0 
    input [9:0] Pix_406, // sfix10_En0 
    input [9:0] Pix_407, // sfix10_En0 
    input [9:0] Pix_408, // sfix10_En0 
    input [9:0] Pix_409, // sfix10_En0 
    input [9:0] Pix_410, // sfix10_En0 
    input [9:0] Pix_411, // sfix10_En0 
    input [9:0] Pix_412, // sfix10_En0 
    input [9:0] Pix_413, // sfix10_En0 
    input [9:0] Pix_414, // sfix10_En0 
    input [9:0] Pix_415, // sfix10_En0 
    input [9:0] Pix_416, // sfix10_En0 
    input [9:0] Pix_417, // sfix10_En0 
    input [9:0] Pix_418, // sfix10_En0 
    input [9:0] Pix_419, // sfix10_En0 
    input [9:0] Pix_420, // sfix10_En0 
    input [9:0] Pix_421, // sfix10_En0 
    input [9:0] Pix_422, // sfix10_En0 
    input [9:0] Pix_423, // sfix10_En0 
    input [9:0] Pix_424, // sfix10_En0 
    input [9:0] Pix_425, // sfix10_En0 
    input [9:0] Pix_426, // sfix10_En0 
    input [9:0] Pix_427, // sfix10_En0 
    input [9:0] Pix_428, // sfix10_En0 
    input [9:0] Pix_429, // sfix10_En0 
    input [9:0] Pix_430, // sfix10_En0 
    input [9:0] Pix_431, // sfix10_En0 
    input [9:0] Pix_432, // sfix10_En0 
    input [9:0] Pix_433, // sfix10_En0 
    input [9:0] Pix_434, // sfix10_En0 
    input [9:0] Pix_435, // sfix10_En0 
    input [9:0] Pix_436, // sfix10_En0 
    input [9:0] Pix_437, // sfix10_En0 
    input [9:0] Pix_438, // sfix10_En0 
    input [9:0] Pix_439, // sfix10_En0 
    input [9:0] Pix_440, // sfix10_En0 
    input [9:0] Pix_441, // sfix10_En0 
    input [9:0] Pix_442, // sfix10_En0 
    input [9:0] Pix_443, // sfix10_En0 
    input [9:0] Pix_444, // sfix10_En0 
    input [9:0] Pix_445, // sfix10_En0 
    input [9:0] Pix_446, // sfix10_En0 
    input [9:0] Pix_447, // sfix10_En0 
    input [9:0] Pix_448, // sfix10_En0 
    input [9:0] Pix_449, // sfix10_En0 
    input [9:0] Pix_450, // sfix10_En0 
    input [9:0] Pix_451, // sfix10_En0 
    input [9:0] Pix_452, // sfix10_En0 
    input [9:0] Pix_453, // sfix10_En0 
    input [9:0] Pix_454, // sfix10_En0 
    input [9:0] Pix_455, // sfix10_En0 
    input [9:0] Pix_456, // sfix10_En0 
    input [9:0] Pix_457, // sfix10_En0 
    input [9:0] Pix_458, // sfix10_En0 
    input [9:0] Pix_459, // sfix10_En0 
    input [9:0] Pix_460, // sfix10_En0 
    input [9:0] Pix_461, // sfix10_En0 
    input [9:0] Pix_462, // sfix10_En0 
    input [9:0] Pix_463, // sfix10_En0 
    input [9:0] Pix_464, // sfix10_En0 
    input [9:0] Pix_465, // sfix10_En0 
    input [9:0] Pix_466, // sfix10_En0 
    input [9:0] Pix_467, // sfix10_En0 
    input [9:0] Pix_468, // sfix10_En0 
    input [9:0] Pix_469, // sfix10_En0 
    input [9:0] Pix_470, // sfix10_En0 
    input [9:0] Pix_471, // sfix10_En0 
    input [9:0] Pix_472, // sfix10_En0 
    input [9:0] Pix_473, // sfix10_En0 
    input [9:0] Pix_474, // sfix10_En0 
    input [9:0] Pix_475, // sfix10_En0 
    input [9:0] Pix_476, // sfix10_En0 
    input [9:0] Pix_477, // sfix10_En0 
    input [9:0] Pix_478, // sfix10_En0 
    input [9:0] Pix_479, // sfix10_En0 
    input [9:0] Pix_480, // sfix10_En0 
    input [9:0] Pix_481, // sfix10_En0 
    input [9:0] Pix_482, // sfix10_En0 
    input [9:0] Pix_483, // sfix10_En0 
    input [9:0] Pix_484, // sfix10_En0 
    input [9:0] Pix_485, // sfix10_En0 
    input [9:0] Pix_486, // sfix10_En0 
    input [9:0] Pix_487, // sfix10_En0 
    input [9:0] Pix_488, // sfix10_En0 
    input [9:0] Pix_489, // sfix10_En0 
    input [9:0] Pix_490, // sfix10_En0 
    input [9:0] Pix_491, // sfix10_En0 
    input [9:0] Pix_492, // sfix10_En0 
    input [9:0] Pix_493, // sfix10_En0 
    input [9:0] Pix_494, // sfix10_En0 
    input [9:0] Pix_495, // sfix10_En0 
    input [9:0] Pix_496, // sfix10_En0 
    input [9:0] Pix_497, // sfix10_En0 
    input [9:0] Pix_498, // sfix10_En0 
    input [9:0] Pix_499, // sfix10_En0 
    input [9:0] Pix_500, // sfix10_En0 
    input [9:0] Pix_501, // sfix10_En0 
    input [9:0] Pix_502, // sfix10_En0 
    input [9:0] Pix_503, // sfix10_En0 
    input [9:0] Pix_504, // sfix10_En0 
    input [9:0] Pix_505, // sfix10_En0 
    input [9:0] Pix_506, // sfix10_En0 
    input [9:0] Pix_507, // sfix10_En0 
    input [9:0] Pix_508, // sfix10_En0 
    input [9:0] Pix_509, // sfix10_En0 
    input [9:0] Pix_510, // sfix10_En0 
    input [9:0] Pix_511, // sfix10_En0 
    input [9:0] Pix_512, // sfix10_En0 
    input [9:0] Pix_513, // sfix10_En0 
    input [9:0] Pix_514, // sfix10_En0 
    input [9:0] Pix_515, // sfix10_En0 
    input [9:0] Pix_516, // sfix10_En0 
    input [9:0] Pix_517, // sfix10_En0 
    input [9:0] Pix_518, // sfix10_En0 
    input [9:0] Pix_519, // sfix10_En0 
    input [9:0] Pix_520, // sfix10_En0 
    input [9:0] Pix_521, // sfix10_En0 
    input [9:0] Pix_522, // sfix10_En0 
    input [9:0] Pix_523, // sfix10_En0 
    input [9:0] Pix_524, // sfix10_En0 
    input [9:0] Pix_525, // sfix10_En0 
    input [9:0] Pix_526, // sfix10_En0 
    input [9:0] Pix_527, // sfix10_En0 
    input [9:0] Pix_528, // sfix10_En0 
    input [9:0] Pix_529, // sfix10_En0 
    input [9:0] Pix_530, // sfix10_En0 
    input [9:0] Pix_531, // sfix10_En0 
    input [9:0] Pix_532, // sfix10_En0 
    input [9:0] Pix_533, // sfix10_En0 
    input [9:0] Pix_534, // sfix10_En0 
    input [9:0] Pix_535, // sfix10_En0 
    input [9:0] Pix_536, // sfix10_En0 
    input [9:0] Pix_537, // sfix10_En0 
    input [9:0] Pix_538, // sfix10_En0 
    input [9:0] Pix_539, // sfix10_En0 
    input [9:0] Pix_540, // sfix10_En0 
    input [9:0] Pix_541, // sfix10_En0 
    input [9:0] Pix_542, // sfix10_En0 
    input [9:0] Pix_543, // sfix10_En0 
    input [9:0] Pix_544, // sfix10_En0 
    input [9:0] Pix_545, // sfix10_En0 
    input [9:0] Pix_546, // sfix10_En0 
    input [9:0] Pix_547, // sfix10_En0 
    input [9:0] Pix_548, // sfix10_En0 
    input [9:0] Pix_549, // sfix10_En0 
    input [9:0] Pix_550, // sfix10_En0 
    input [9:0] Pix_551, // sfix10_En0 
    input [9:0] Pix_552, // sfix10_En0 
    input [9:0] Pix_553, // sfix10_En0 
    input [9:0] Pix_554, // sfix10_En0 
    input [9:0] Pix_555, // sfix10_En0 
    input [9:0] Pix_556, // sfix10_En0 
    input [9:0] Pix_557, // sfix10_En0 
    input [9:0] Pix_558, // sfix10_En0 
    input [9:0] Pix_559, // sfix10_En0 
    input [9:0] Pix_560, // sfix10_En0 
    input [9:0] Pix_561, // sfix10_En0 
    input [9:0] Pix_562, // sfix10_En0 
    input [9:0] Pix_563, // sfix10_En0 
    input [9:0] Pix_564, // sfix10_En0 
    input [9:0] Pix_565, // sfix10_En0 
    input [9:0] Pix_566, // sfix10_En0 
    input [9:0] Pix_567, // sfix10_En0 
    input [9:0] Pix_568, // sfix10_En0 
    input [9:0] Pix_569, // sfix10_En0 
    input [9:0] Pix_570, // sfix10_En0 
    input [9:0] Pix_571, // sfix10_En0 
    input [9:0] Pix_572, // sfix10_En0 
    input [9:0] Pix_573, // sfix10_En0 
    input [9:0] Pix_574, // sfix10_En0 
    input [9:0] Pix_575, // sfix10_En0 
    input [9:0] Pix_576, // sfix10_En0 
    input [9:0] Pix_577, // sfix10_En0 
    input [9:0] Pix_578, // sfix10_En0 
    input [9:0] Pix_579, // sfix10_En0 
    input [9:0] Pix_580, // sfix10_En0 
    input [9:0] Pix_581, // sfix10_En0 
    input [9:0] Pix_582, // sfix10_En0 
    input [9:0] Pix_583, // sfix10_En0 
    input [9:0] Pix_584, // sfix10_En0 
    input [9:0] Pix_585, // sfix10_En0 
    input [9:0] Pix_586, // sfix10_En0 
    input [9:0] Pix_587, // sfix10_En0 
    input [9:0] Pix_588, // sfix10_En0 
    input [9:0] Pix_589, // sfix10_En0 
    input [9:0] Pix_590, // sfix10_En0 
    input [9:0] Pix_591, // sfix10_En0 
    input [9:0] Pix_592, // sfix10_En0 
    input [9:0] Pix_593, // sfix10_En0 
    input [9:0] Pix_594, // sfix10_En0 
    input [9:0] Pix_595, // sfix10_En0 
    input [9:0] Pix_596, // sfix10_En0 
    input [9:0] Pix_597, // sfix10_En0 
    input [9:0] Pix_598, // sfix10_En0 
    input [9:0] Pix_599, // sfix10_En0 
    input [9:0] Pix_600, // sfix10_En0 
    input [9:0] Pix_601, // sfix10_En0 
    input [9:0] Pix_602, // sfix10_En0 
    input [9:0] Pix_603, // sfix10_En0 
    input [9:0] Pix_604, // sfix10_En0 
    input [9:0] Pix_605, // sfix10_En0 
    input [9:0] Pix_606, // sfix10_En0 
    input [9:0] Pix_607, // sfix10_En0 
    input [9:0] Pix_608, // sfix10_En0 
    input [9:0] Pix_609, // sfix10_En0 
    input [9:0] Pix_610, // sfix10_En0 
    input [9:0] Pix_611, // sfix10_En0 
    input [9:0] Pix_612, // sfix10_En0 
    input [9:0] Pix_613, // sfix10_En0 
    input [9:0] Pix_614, // sfix10_En0 
    input [9:0] Pix_615, // sfix10_En0 
    input [9:0] Pix_616, // sfix10_En0 
    input [9:0] Pix_617, // sfix10_En0 
    input [9:0] Pix_618, // sfix10_En0 
    input [9:0] Pix_619, // sfix10_En0 
    input [9:0] Pix_620, // sfix10_En0 
    input [9:0] Pix_621, // sfix10_En0 
    input [9:0] Pix_622, // sfix10_En0 
    input [9:0] Pix_623, // sfix10_En0 
    input [9:0] Pix_624, // sfix10_En0 
    input [9:0] Pix_625, // sfix10_En0 
    input [9:0] Pix_626, // sfix10_En0 
    input [9:0] Pix_627, // sfix10_En0 
    input [9:0] Pix_628, // sfix10_En0 
    input [9:0] Pix_629, // sfix10_En0 
    input [9:0] Pix_630, // sfix10_En0 
    input [9:0] Pix_631, // sfix10_En0 
    input [9:0] Pix_632, // sfix10_En0 
    input [9:0] Pix_633, // sfix10_En0 
    input [9:0] Pix_634, // sfix10_En0 
    input [9:0] Pix_635, // sfix10_En0 
    input [9:0] Pix_636, // sfix10_En0 
    input [9:0] Pix_637, // sfix10_En0 
    input [9:0] Pix_638, // sfix10_En0 
    input [9:0] Pix_639, // sfix10_En0 
    input [9:0] Pix_640, // sfix10_En0 
    input [9:0] Pix_641, // sfix10_En0 
    input [9:0] Pix_642, // sfix10_En0 
    input [9:0] Pix_643, // sfix10_En0 
    input [9:0] Pix_644, // sfix10_En0 
    input [9:0] Pix_645, // sfix10_En0 
    input [9:0] Pix_646, // sfix10_En0 
    input [9:0] Pix_647, // sfix10_En0 
    input [9:0] Pix_648, // sfix10_En0 
    input [9:0] Pix_649, // sfix10_En0 
    input [9:0] Pix_650, // sfix10_En0 
    input [9:0] Pix_651, // sfix10_En0 
    input [9:0] Pix_652, // sfix10_En0 
    input [9:0] Pix_653, // sfix10_En0 
    input [9:0] Pix_654, // sfix10_En0 
    input [9:0] Pix_655, // sfix10_En0 
    input [9:0] Pix_656, // sfix10_En0 
    input [9:0] Pix_657, // sfix10_En0 
    input [9:0] Pix_658, // sfix10_En0 
    input [9:0] Pix_659, // sfix10_En0 
    input [9:0] Pix_660, // sfix10_En0 
    input [9:0] Pix_661, // sfix10_En0 
    input [9:0] Pix_662, // sfix10_En0 
    input [9:0] Pix_663, // sfix10_En0 
    input [9:0] Pix_664, // sfix10_En0 
    input [9:0] Pix_665, // sfix10_En0 
    input [9:0] Pix_666, // sfix10_En0 
    input [9:0] Pix_667, // sfix10_En0 
    input [9:0] Pix_668, // sfix10_En0 
    input [9:0] Pix_669, // sfix10_En0 
    input [9:0] Pix_670, // sfix10_En0 
    input [9:0] Pix_671, // sfix10_En0 
    input [9:0] Pix_672, // sfix10_En0 
    input [9:0] Pix_673, // sfix10_En0 
    input [9:0] Pix_674, // sfix10_En0 
    input [9:0] Pix_675, // sfix10_En0 
    input [9:0] Pix_676, // sfix10_En0 
    input [9:0] Pix_677, // sfix10_En0 
    input [9:0] Pix_678, // sfix10_En0 
    input [9:0] Pix_679, // sfix10_En0 
    input [9:0] Pix_680, // sfix10_En0 
    input [9:0] Pix_681, // sfix10_En0 
    input [9:0] Pix_682, // sfix10_En0 
    input [9:0] Pix_683, // sfix10_En0 
    input [9:0] Pix_684, // sfix10_En0 
    input [9:0] Pix_685, // sfix10_En0 
    input [9:0] Pix_686, // sfix10_En0 
    input [9:0] Pix_687, // sfix10_En0 
    input [9:0] Pix_688, // sfix10_En0 
    input [9:0] Pix_689, // sfix10_En0 
    input [9:0] Pix_690, // sfix10_En0 
    input [9:0] Pix_691, // sfix10_En0 
    input [9:0] Pix_692, // sfix10_En0 
    input [9:0] Pix_693, // sfix10_En0 
    input [9:0] Pix_694, // sfix10_En0 
    input [9:0] Pix_695, // sfix10_En0 
    input [9:0] Pix_696, // sfix10_En0 
    input [9:0] Pix_697, // sfix10_En0 
    input [9:0] Pix_698, // sfix10_En0 
    input [9:0] Pix_699, // sfix10_En0 
    input [9:0] Pix_700, // sfix10_En0 
    input [9:0] Pix_701, // sfix10_En0 
    input [9:0] Pix_702, // sfix10_En0 
    input [9:0] Pix_703, // sfix10_En0 
    input [9:0] Pix_704, // sfix10_En0 
    input [9:0] Pix_705, // sfix10_En0 
    input [9:0] Pix_706, // sfix10_En0 
    input [9:0] Pix_707, // sfix10_En0 
    input [9:0] Pix_708, // sfix10_En0 
    input [9:0] Pix_709, // sfix10_En0 
    input [9:0] Pix_710, // sfix10_En0 
    input [9:0] Pix_711, // sfix10_En0 
    input [9:0] Pix_712, // sfix10_En0 
    input [9:0] Pix_713, // sfix10_En0 
    input [9:0] Pix_714, // sfix10_En0 
    input [9:0] Pix_715, // sfix10_En0 
    input [9:0] Pix_716, // sfix10_En0 
    input [9:0] Pix_717, // sfix10_En0 
    input [9:0] Pix_718, // sfix10_En0 
    input [9:0] Pix_719, // sfix10_En0 
    input [9:0] Pix_720, // sfix10_En0 
    input [9:0] Pix_721, // sfix10_En0 
    input [9:0] Pix_722, // sfix10_En0 
    input [9:0] Pix_723, // sfix10_En0 
    input [9:0] Pix_724, // sfix10_En0 
    input [9:0] Pix_725, // sfix10_En0 
    input [9:0] Pix_726, // sfix10_En0 
    input [9:0] Pix_727, // sfix10_En0 
    input [9:0] Pix_728, // sfix10_En0 
    input [9:0] Pix_729, // sfix10_En0 
    input [9:0] Pix_730, // sfix10_En0 
    input [9:0] Pix_731, // sfix10_En0 
    input [9:0] Pix_732, // sfix10_En0 
    input [9:0] Pix_733, // sfix10_En0 
    input [9:0] Pix_734, // sfix10_En0 
    input [9:0] Pix_735, // sfix10_En0 
    input [9:0] Pix_736, // sfix10_En0 
    input [9:0] Pix_737, // sfix10_En0 
    input [9:0] Pix_738, // sfix10_En0 
    input [9:0] Pix_739, // sfix10_En0 
    input [9:0] Pix_740, // sfix10_En0 
    input [9:0] Pix_741, // sfix10_En0 
    input [9:0] Pix_742, // sfix10_En0 
    input [9:0] Pix_743, // sfix10_En0 
    input [9:0] Pix_744, // sfix10_En0 
    input [9:0] Pix_745, // sfix10_En0 
    input [9:0] Pix_746, // sfix10_En0 
    input [9:0] Pix_747, // sfix10_En0 
    input [9:0] Pix_748, // sfix10_En0 
    input [9:0] Pix_749, // sfix10_En0 
    input [9:0] Pix_750, // sfix10_En0 
    input [9:0] Pix_751, // sfix10_En0 
    input [9:0] Pix_752, // sfix10_En0 
    input [9:0] Pix_753, // sfix10_En0 
    input [9:0] Pix_754, // sfix10_En0 
    input [9:0] Pix_755, // sfix10_En0 
    input [9:0] Pix_756, // sfix10_En0 
    input [9:0] Pix_757, // sfix10_En0 
    input [9:0] Pix_758, // sfix10_En0 
    input [9:0] Pix_759, // sfix10_En0 
    input [9:0] Pix_760, // sfix10_En0 
    input [9:0] Pix_761, // sfix10_En0 
    input [9:0] Pix_762, // sfix10_En0 
    input [9:0] Pix_763, // sfix10_En0 
    input [9:0] Pix_764, // sfix10_En0 
    input [9:0] Pix_765, // sfix10_En0 
    input [9:0] Pix_766, // sfix10_En0 
    input [9:0] Pix_767, // sfix10_En0 
    input [9:0] Pix_768, // sfix10_En0 
    input [9:0] Pix_769, // sfix10_En0 
    input [9:0] Pix_770, // sfix10_En0 
    input [9:0] Pix_771, // sfix10_En0 
    input [9:0] Pix_772, // sfix10_En0 
    input [9:0] Pix_773, // sfix10_En0 
    input [9:0] Pix_774, // sfix10_En0 
    input [9:0] Pix_775, // sfix10_En0 
    input [9:0] Pix_776, // sfix10_En0 
    input [9:0] Pix_777, // sfix10_En0 
    input [9:0] Pix_778, // sfix10_En0 
    input [9:0] Pix_779, // sfix10_En0 
    input [9:0] Pix_780, // sfix10_En0 
    input [9:0] Pix_781, // sfix10_En0 
    input [9:0] Pix_782, // sfix10_En0 
    input [9:0] Pix_783, // sfix10_En0 
    input [9:0] Pix_784, // sfix10_En0 ?
    output [3:0] Image_Number, // sfix26_En18 
    output Output_Valid 
 );

// active low reset 
wire GlobalResetn = ~GlobalReset;

// buffered image
reg [`PIX_WIDTH-1:0] Pixels [0:784];

// initialize pixels when Input_Valid 0 --> 1
always @ (posedge Input_Valid) begin
    Pixels[0] <= Pix_0[`PIX_WIDTH-1:0];
    Pixels[1] <= Pix_1[`PIX_WIDTH-1:0];
    Pixels[2] <= Pix_2[`PIX_WIDTH-1:0];
    Pixels[3] <= Pix_3[`PIX_WIDTH-1:0];
    Pixels[4] <= Pix_4[`PIX_WIDTH-1:0];
    Pixels[5] <= Pix_5[`PIX_WIDTH-1:0];
    Pixels[6] <= Pix_6[`PIX_WIDTH-1:0];
    Pixels[7] <= Pix_7[`PIX_WIDTH-1:0];
    Pixels[8] <= Pix_8[`PIX_WIDTH-1:0];
    Pixels[9] <= Pix_9[`PIX_WIDTH-1:0];
    Pixels[10] <= Pix_10[`PIX_WIDTH-1:0];
    Pixels[11] <= Pix_11[`PIX_WIDTH-1:0];
    Pixels[12] <= Pix_12[`PIX_WIDTH-1:0];
    Pixels[13] <= Pix_13[`PIX_WIDTH-1:0];
    Pixels[14] <= Pix_14[`PIX_WIDTH-1:0];
    Pixels[15] <= Pix_15[`PIX_WIDTH-1:0];
    Pixels[16] <= Pix_16[`PIX_WIDTH-1:0];
    Pixels[17] <= Pix_17[`PIX_WIDTH-1:0];
    Pixels[18] <= Pix_18[`PIX_WIDTH-1:0];
    Pixels[19] <= Pix_19[`PIX_WIDTH-1:0];
    Pixels[20] <= Pix_20[`PIX_WIDTH-1:0];
    Pixels[21] <= Pix_21[`PIX_WIDTH-1:0];
    Pixels[22] <= Pix_22[`PIX_WIDTH-1:0];
    Pixels[23] <= Pix_23[`PIX_WIDTH-1:0];
    Pixels[24] <= Pix_24[`PIX_WIDTH-1:0];
    Pixels[25] <= Pix_25[`PIX_WIDTH-1:0];
    Pixels[26] <= Pix_26[`PIX_WIDTH-1:0];
    Pixels[27] <= Pix_27[`PIX_WIDTH-1:0];
    Pixels[28] <= Pix_28[`PIX_WIDTH-1:0];
    Pixels[29] <= Pix_29[`PIX_WIDTH-1:0];
    Pixels[30] <= Pix_30[`PIX_WIDTH-1:0];
    Pixels[31] <= Pix_31[`PIX_WIDTH-1:0];
    Pixels[32] <= Pix_32[`PIX_WIDTH-1:0];
    Pixels[33] <= Pix_33[`PIX_WIDTH-1:0];
    Pixels[34] <= Pix_34[`PIX_WIDTH-1:0];
    Pixels[35] <= Pix_35[`PIX_WIDTH-1:0];
    Pixels[36] <= Pix_36[`PIX_WIDTH-1:0];
    Pixels[37] <= Pix_37[`PIX_WIDTH-1:0];
    Pixels[38] <= Pix_38[`PIX_WIDTH-1:0];
    Pixels[39] <= Pix_39[`PIX_WIDTH-1:0];
    Pixels[40] <= Pix_40[`PIX_WIDTH-1:0];
    Pixels[41] <= Pix_41[`PIX_WIDTH-1:0];
    Pixels[42] <= Pix_42[`PIX_WIDTH-1:0];
    Pixels[43] <= Pix_43[`PIX_WIDTH-1:0];
    Pixels[44] <= Pix_44[`PIX_WIDTH-1:0];
    Pixels[45] <= Pix_45[`PIX_WIDTH-1:0];
    Pixels[46] <= Pix_46[`PIX_WIDTH-1:0];
    Pixels[47] <= Pix_47[`PIX_WIDTH-1:0];
    Pixels[48] <= Pix_48[`PIX_WIDTH-1:0];
    Pixels[49] <= Pix_49[`PIX_WIDTH-1:0];
    Pixels[50] <= Pix_50[`PIX_WIDTH-1:0];
    Pixels[51] <= Pix_51[`PIX_WIDTH-1:0];
    Pixels[52] <= Pix_52[`PIX_WIDTH-1:0];
    Pixels[53] <= Pix_53[`PIX_WIDTH-1:0];
    Pixels[54] <= Pix_54[`PIX_WIDTH-1:0];
    Pixels[55] <= Pix_55[`PIX_WIDTH-1:0];
    Pixels[56] <= Pix_56[`PIX_WIDTH-1:0];
    Pixels[57] <= Pix_57[`PIX_WIDTH-1:0];
    Pixels[58] <= Pix_58[`PIX_WIDTH-1:0];
    Pixels[59] <= Pix_59[`PIX_WIDTH-1:0];
    Pixels[60] <= Pix_60[`PIX_WIDTH-1:0];
    Pixels[61] <= Pix_61[`PIX_WIDTH-1:0];
    Pixels[62] <= Pix_62[`PIX_WIDTH-1:0];
    Pixels[63] <= Pix_63[`PIX_WIDTH-1:0];
    Pixels[64] <= Pix_64[`PIX_WIDTH-1:0];
    Pixels[65] <= Pix_65[`PIX_WIDTH-1:0];
    Pixels[66] <= Pix_66[`PIX_WIDTH-1:0];
    Pixels[67] <= Pix_67[`PIX_WIDTH-1:0];
    Pixels[68] <= Pix_68[`PIX_WIDTH-1:0];
    Pixels[69] <= Pix_69[`PIX_WIDTH-1:0];
    Pixels[70] <= Pix_70[`PIX_WIDTH-1:0];
    Pixels[71] <= Pix_71[`PIX_WIDTH-1:0];
    Pixels[72] <= Pix_72[`PIX_WIDTH-1:0];
    Pixels[73] <= Pix_73[`PIX_WIDTH-1:0];
    Pixels[74] <= Pix_74[`PIX_WIDTH-1:0];
    Pixels[75] <= Pix_75[`PIX_WIDTH-1:0];
    Pixels[76] <= Pix_76[`PIX_WIDTH-1:0];
    Pixels[77] <= Pix_77[`PIX_WIDTH-1:0];
    Pixels[78] <= Pix_78[`PIX_WIDTH-1:0];
    Pixels[79] <= Pix_79[`PIX_WIDTH-1:0];
    Pixels[80] <= Pix_80[`PIX_WIDTH-1:0];
    Pixels[81] <= Pix_81[`PIX_WIDTH-1:0];
    Pixels[82] <= Pix_82[`PIX_WIDTH-1:0];
    Pixels[83] <= Pix_83[`PIX_WIDTH-1:0];
    Pixels[84] <= Pix_84[`PIX_WIDTH-1:0];
    Pixels[85] <= Pix_85[`PIX_WIDTH-1:0];
    Pixels[86] <= Pix_86[`PIX_WIDTH-1:0];
    Pixels[87] <= Pix_87[`PIX_WIDTH-1:0];
    Pixels[88] <= Pix_88[`PIX_WIDTH-1:0];
    Pixels[89] <= Pix_89[`PIX_WIDTH-1:0];
    Pixels[90] <= Pix_90[`PIX_WIDTH-1:0];
    Pixels[91] <= Pix_91[`PIX_WIDTH-1:0];
    Pixels[92] <= Pix_92[`PIX_WIDTH-1:0];
    Pixels[93] <= Pix_93[`PIX_WIDTH-1:0];
    Pixels[94] <= Pix_94[`PIX_WIDTH-1:0];
    Pixels[95] <= Pix_95[`PIX_WIDTH-1:0];
    Pixels[96] <= Pix_96[`PIX_WIDTH-1:0];
    Pixels[97] <= Pix_97[`PIX_WIDTH-1:0];
    Pixels[98] <= Pix_98[`PIX_WIDTH-1:0];
    Pixels[99] <= Pix_99[`PIX_WIDTH-1:0];
    Pixels[100] <= Pix_100[`PIX_WIDTH-1:0];
    Pixels[101] <= Pix_101[`PIX_WIDTH-1:0];
    Pixels[102] <= Pix_102[`PIX_WIDTH-1:0];
    Pixels[103] <= Pix_103[`PIX_WIDTH-1:0];
    Pixels[104] <= Pix_104[`PIX_WIDTH-1:0];
    Pixels[105] <= Pix_105[`PIX_WIDTH-1:0];
    Pixels[106] <= Pix_106[`PIX_WIDTH-1:0];
    Pixels[107] <= Pix_107[`PIX_WIDTH-1:0];
    Pixels[108] <= Pix_108[`PIX_WIDTH-1:0];
    Pixels[109] <= Pix_109[`PIX_WIDTH-1:0];
    Pixels[110] <= Pix_110[`PIX_WIDTH-1:0];
    Pixels[111] <= Pix_111[`PIX_WIDTH-1:0];
    Pixels[112] <= Pix_112[`PIX_WIDTH-1:0];
    Pixels[113] <= Pix_113[`PIX_WIDTH-1:0];
    Pixels[114] <= Pix_114[`PIX_WIDTH-1:0];
    Pixels[115] <= Pix_115[`PIX_WIDTH-1:0];
    Pixels[116] <= Pix_116[`PIX_WIDTH-1:0];
    Pixels[117] <= Pix_117[`PIX_WIDTH-1:0];
    Pixels[118] <= Pix_118[`PIX_WIDTH-1:0];
    Pixels[119] <= Pix_119[`PIX_WIDTH-1:0];
    Pixels[120] <= Pix_120[`PIX_WIDTH-1:0];
    Pixels[121] <= Pix_121[`PIX_WIDTH-1:0];
    Pixels[122] <= Pix_122[`PIX_WIDTH-1:0];
    Pixels[123] <= Pix_123[`PIX_WIDTH-1:0];
    Pixels[124] <= Pix_124[`PIX_WIDTH-1:0];
    Pixels[125] <= Pix_125[`PIX_WIDTH-1:0];
    Pixels[126] <= Pix_126[`PIX_WIDTH-1:0];
    Pixels[127] <= Pix_127[`PIX_WIDTH-1:0];
    Pixels[128] <= Pix_128[`PIX_WIDTH-1:0];
    Pixels[129] <= Pix_129[`PIX_WIDTH-1:0];
    Pixels[130] <= Pix_130[`PIX_WIDTH-1:0];
    Pixels[131] <= Pix_131[`PIX_WIDTH-1:0];
    Pixels[132] <= Pix_132[`PIX_WIDTH-1:0];
    Pixels[133] <= Pix_133[`PIX_WIDTH-1:0];
    Pixels[134] <= Pix_134[`PIX_WIDTH-1:0];
    Pixels[135] <= Pix_135[`PIX_WIDTH-1:0];
    Pixels[136] <= Pix_136[`PIX_WIDTH-1:0];
    Pixels[137] <= Pix_137[`PIX_WIDTH-1:0];
    Pixels[138] <= Pix_138[`PIX_WIDTH-1:0];
    Pixels[139] <= Pix_139[`PIX_WIDTH-1:0];
    Pixels[140] <= Pix_140[`PIX_WIDTH-1:0];
    Pixels[141] <= Pix_141[`PIX_WIDTH-1:0];
    Pixels[142] <= Pix_142[`PIX_WIDTH-1:0];
    Pixels[143] <= Pix_143[`PIX_WIDTH-1:0];
    Pixels[144] <= Pix_144[`PIX_WIDTH-1:0];
    Pixels[145] <= Pix_145[`PIX_WIDTH-1:0];
    Pixels[146] <= Pix_146[`PIX_WIDTH-1:0];
    Pixels[147] <= Pix_147[`PIX_WIDTH-1:0];
    Pixels[148] <= Pix_148[`PIX_WIDTH-1:0];
    Pixels[149] <= Pix_149[`PIX_WIDTH-1:0];
    Pixels[150] <= Pix_150[`PIX_WIDTH-1:0];
    Pixels[151] <= Pix_151[`PIX_WIDTH-1:0];
    Pixels[152] <= Pix_152[`PIX_WIDTH-1:0];
    Pixels[153] <= Pix_153[`PIX_WIDTH-1:0];
    Pixels[154] <= Pix_154[`PIX_WIDTH-1:0];
    Pixels[155] <= Pix_155[`PIX_WIDTH-1:0];
    Pixels[156] <= Pix_156[`PIX_WIDTH-1:0];
    Pixels[157] <= Pix_157[`PIX_WIDTH-1:0];
    Pixels[158] <= Pix_158[`PIX_WIDTH-1:0];
    Pixels[159] <= Pix_159[`PIX_WIDTH-1:0];
    Pixels[160] <= Pix_160[`PIX_WIDTH-1:0];
    Pixels[161] <= Pix_161[`PIX_WIDTH-1:0];
    Pixels[162] <= Pix_162[`PIX_WIDTH-1:0];
    Pixels[163] <= Pix_163[`PIX_WIDTH-1:0];
    Pixels[164] <= Pix_164[`PIX_WIDTH-1:0];
    Pixels[165] <= Pix_165[`PIX_WIDTH-1:0];
    Pixels[166] <= Pix_166[`PIX_WIDTH-1:0];
    Pixels[167] <= Pix_167[`PIX_WIDTH-1:0];
    Pixels[168] <= Pix_168[`PIX_WIDTH-1:0];
    Pixels[169] <= Pix_169[`PIX_WIDTH-1:0];
    Pixels[170] <= Pix_170[`PIX_WIDTH-1:0];
    Pixels[171] <= Pix_171[`PIX_WIDTH-1:0];
    Pixels[172] <= Pix_172[`PIX_WIDTH-1:0];
    Pixels[173] <= Pix_173[`PIX_WIDTH-1:0];
    Pixels[174] <= Pix_174[`PIX_WIDTH-1:0];
    Pixels[175] <= Pix_175[`PIX_WIDTH-1:0];
    Pixels[176] <= Pix_176[`PIX_WIDTH-1:0];
    Pixels[177] <= Pix_177[`PIX_WIDTH-1:0];
    Pixels[178] <= Pix_178[`PIX_WIDTH-1:0];
    Pixels[179] <= Pix_179[`PIX_WIDTH-1:0];
    Pixels[180] <= Pix_180[`PIX_WIDTH-1:0];
    Pixels[181] <= Pix_181[`PIX_WIDTH-1:0];
    Pixels[182] <= Pix_182[`PIX_WIDTH-1:0];
    Pixels[183] <= Pix_183[`PIX_WIDTH-1:0];
    Pixels[184] <= Pix_184[`PIX_WIDTH-1:0];
    Pixels[185] <= Pix_185[`PIX_WIDTH-1:0];
    Pixels[186] <= Pix_186[`PIX_WIDTH-1:0];
    Pixels[187] <= Pix_187[`PIX_WIDTH-1:0];
    Pixels[188] <= Pix_188[`PIX_WIDTH-1:0];
    Pixels[189] <= Pix_189[`PIX_WIDTH-1:0];
    Pixels[190] <= Pix_190[`PIX_WIDTH-1:0];
    Pixels[191] <= Pix_191[`PIX_WIDTH-1:0];
    Pixels[192] <= Pix_192[`PIX_WIDTH-1:0];
    Pixels[193] <= Pix_193[`PIX_WIDTH-1:0];
    Pixels[194] <= Pix_194[`PIX_WIDTH-1:0];
    Pixels[195] <= Pix_195[`PIX_WIDTH-1:0];
    Pixels[196] <= Pix_196[`PIX_WIDTH-1:0];
    Pixels[197] <= Pix_197[`PIX_WIDTH-1:0];
    Pixels[198] <= Pix_198[`PIX_WIDTH-1:0];
    Pixels[199] <= Pix_199[`PIX_WIDTH-1:0];
    Pixels[200] <= Pix_200[`PIX_WIDTH-1:0];
    Pixels[201] <= Pix_201[`PIX_WIDTH-1:0];
    Pixels[202] <= Pix_202[`PIX_WIDTH-1:0];
    Pixels[203] <= Pix_203[`PIX_WIDTH-1:0];
    Pixels[204] <= Pix_204[`PIX_WIDTH-1:0];
    Pixels[205] <= Pix_205[`PIX_WIDTH-1:0];
    Pixels[206] <= Pix_206[`PIX_WIDTH-1:0];
    Pixels[207] <= Pix_207[`PIX_WIDTH-1:0];
    Pixels[208] <= Pix_208[`PIX_WIDTH-1:0];
    Pixels[209] <= Pix_209[`PIX_WIDTH-1:0];
    Pixels[210] <= Pix_210[`PIX_WIDTH-1:0];
    Pixels[211] <= Pix_211[`PIX_WIDTH-1:0];
    Pixels[212] <= Pix_212[`PIX_WIDTH-1:0];
    Pixels[213] <= Pix_213[`PIX_WIDTH-1:0];
    Pixels[214] <= Pix_214[`PIX_WIDTH-1:0];
    Pixels[215] <= Pix_215[`PIX_WIDTH-1:0];
    Pixels[216] <= Pix_216[`PIX_WIDTH-1:0];
    Pixels[217] <= Pix_217[`PIX_WIDTH-1:0];
    Pixels[218] <= Pix_218[`PIX_WIDTH-1:0];
    Pixels[219] <= Pix_219[`PIX_WIDTH-1:0];
    Pixels[220] <= Pix_220[`PIX_WIDTH-1:0];
    Pixels[221] <= Pix_221[`PIX_WIDTH-1:0];
    Pixels[222] <= Pix_222[`PIX_WIDTH-1:0];
    Pixels[223] <= Pix_223[`PIX_WIDTH-1:0];
    Pixels[224] <= Pix_224[`PIX_WIDTH-1:0];
    Pixels[225] <= Pix_225[`PIX_WIDTH-1:0];
    Pixels[226] <= Pix_226[`PIX_WIDTH-1:0];
    Pixels[227] <= Pix_227[`PIX_WIDTH-1:0];
    Pixels[228] <= Pix_228[`PIX_WIDTH-1:0];
    Pixels[229] <= Pix_229[`PIX_WIDTH-1:0];
    Pixels[230] <= Pix_230[`PIX_WIDTH-1:0];
    Pixels[231] <= Pix_231[`PIX_WIDTH-1:0];
    Pixels[232] <= Pix_232[`PIX_WIDTH-1:0];
    Pixels[233] <= Pix_233[`PIX_WIDTH-1:0];
    Pixels[234] <= Pix_234[`PIX_WIDTH-1:0];
    Pixels[235] <= Pix_235[`PIX_WIDTH-1:0];
    Pixels[236] <= Pix_236[`PIX_WIDTH-1:0];
    Pixels[237] <= Pix_237[`PIX_WIDTH-1:0];
    Pixels[238] <= Pix_238[`PIX_WIDTH-1:0];
    Pixels[239] <= Pix_239[`PIX_WIDTH-1:0];
    Pixels[240] <= Pix_240[`PIX_WIDTH-1:0];
    Pixels[241] <= Pix_241[`PIX_WIDTH-1:0];
    Pixels[242] <= Pix_242[`PIX_WIDTH-1:0];
    Pixels[243] <= Pix_243[`PIX_WIDTH-1:0];
    Pixels[244] <= Pix_244[`PIX_WIDTH-1:0];
    Pixels[245] <= Pix_245[`PIX_WIDTH-1:0];
    Pixels[246] <= Pix_246[`PIX_WIDTH-1:0];
    Pixels[247] <= Pix_247[`PIX_WIDTH-1:0];
    Pixels[248] <= Pix_248[`PIX_WIDTH-1:0];
    Pixels[249] <= Pix_249[`PIX_WIDTH-1:0];
    Pixels[250] <= Pix_250[`PIX_WIDTH-1:0];
    Pixels[251] <= Pix_251[`PIX_WIDTH-1:0];
    Pixels[252] <= Pix_252[`PIX_WIDTH-1:0];
    Pixels[253] <= Pix_253[`PIX_WIDTH-1:0];
    Pixels[254] <= Pix_254[`PIX_WIDTH-1:0];
    Pixels[255] <= Pix_255[`PIX_WIDTH-1:0];
    Pixels[256] <= Pix_256[`PIX_WIDTH-1:0];
    Pixels[257] <= Pix_257[`PIX_WIDTH-1:0];
    Pixels[258] <= Pix_258[`PIX_WIDTH-1:0];
    Pixels[259] <= Pix_259[`PIX_WIDTH-1:0];
    Pixels[260] <= Pix_260[`PIX_WIDTH-1:0];
    Pixels[261] <= Pix_261[`PIX_WIDTH-1:0];
    Pixels[262] <= Pix_262[`PIX_WIDTH-1:0];
    Pixels[263] <= Pix_263[`PIX_WIDTH-1:0];
    Pixels[264] <= Pix_264[`PIX_WIDTH-1:0];
    Pixels[265] <= Pix_265[`PIX_WIDTH-1:0];
    Pixels[266] <= Pix_266[`PIX_WIDTH-1:0];
    Pixels[267] <= Pix_267[`PIX_WIDTH-1:0];
    Pixels[268] <= Pix_268[`PIX_WIDTH-1:0];
    Pixels[269] <= Pix_269[`PIX_WIDTH-1:0];
    Pixels[270] <= Pix_270[`PIX_WIDTH-1:0];
    Pixels[271] <= Pix_271[`PIX_WIDTH-1:0];
    Pixels[272] <= Pix_272[`PIX_WIDTH-1:0];
    Pixels[273] <= Pix_273[`PIX_WIDTH-1:0];
    Pixels[274] <= Pix_274[`PIX_WIDTH-1:0];
    Pixels[275] <= Pix_275[`PIX_WIDTH-1:0];
    Pixels[276] <= Pix_276[`PIX_WIDTH-1:0];
    Pixels[277] <= Pix_277[`PIX_WIDTH-1:0];
    Pixels[278] <= Pix_278[`PIX_WIDTH-1:0];
    Pixels[279] <= Pix_279[`PIX_WIDTH-1:0];
    Pixels[280] <= Pix_280[`PIX_WIDTH-1:0];
    Pixels[281] <= Pix_281[`PIX_WIDTH-1:0];
    Pixels[282] <= Pix_282[`PIX_WIDTH-1:0];
    Pixels[283] <= Pix_283[`PIX_WIDTH-1:0];
    Pixels[284] <= Pix_284[`PIX_WIDTH-1:0];
    Pixels[285] <= Pix_285[`PIX_WIDTH-1:0];
    Pixels[286] <= Pix_286[`PIX_WIDTH-1:0];
    Pixels[287] <= Pix_287[`PIX_WIDTH-1:0];
    Pixels[288] <= Pix_288[`PIX_WIDTH-1:0];
    Pixels[289] <= Pix_289[`PIX_WIDTH-1:0];
    Pixels[290] <= Pix_290[`PIX_WIDTH-1:0];
    Pixels[291] <= Pix_291[`PIX_WIDTH-1:0];
    Pixels[292] <= Pix_292[`PIX_WIDTH-1:0];
    Pixels[293] <= Pix_293[`PIX_WIDTH-1:0];
    Pixels[294] <= Pix_294[`PIX_WIDTH-1:0];
    Pixels[295] <= Pix_295[`PIX_WIDTH-1:0];
    Pixels[296] <= Pix_296[`PIX_WIDTH-1:0];
    Pixels[297] <= Pix_297[`PIX_WIDTH-1:0];
    Pixels[298] <= Pix_298[`PIX_WIDTH-1:0];
    Pixels[299] <= Pix_299[`PIX_WIDTH-1:0];
    Pixels[300] <= Pix_300[`PIX_WIDTH-1:0];
    Pixels[301] <= Pix_301[`PIX_WIDTH-1:0];
    Pixels[302] <= Pix_302[`PIX_WIDTH-1:0];
    Pixels[303] <= Pix_303[`PIX_WIDTH-1:0];
    Pixels[304] <= Pix_304[`PIX_WIDTH-1:0];
    Pixels[305] <= Pix_305[`PIX_WIDTH-1:0];
    Pixels[306] <= Pix_306[`PIX_WIDTH-1:0];
    Pixels[307] <= Pix_307[`PIX_WIDTH-1:0];
    Pixels[308] <= Pix_308[`PIX_WIDTH-1:0];
    Pixels[309] <= Pix_309[`PIX_WIDTH-1:0];
    Pixels[310] <= Pix_310[`PIX_WIDTH-1:0];
    Pixels[311] <= Pix_311[`PIX_WIDTH-1:0];
    Pixels[312] <= Pix_312[`PIX_WIDTH-1:0];
    Pixels[313] <= Pix_313[`PIX_WIDTH-1:0];
    Pixels[314] <= Pix_314[`PIX_WIDTH-1:0];
    Pixels[315] <= Pix_315[`PIX_WIDTH-1:0];
    Pixels[316] <= Pix_316[`PIX_WIDTH-1:0];
    Pixels[317] <= Pix_317[`PIX_WIDTH-1:0];
    Pixels[318] <= Pix_318[`PIX_WIDTH-1:0];
    Pixels[319] <= Pix_319[`PIX_WIDTH-1:0];
    Pixels[320] <= Pix_320[`PIX_WIDTH-1:0];
    Pixels[321] <= Pix_321[`PIX_WIDTH-1:0];
    Pixels[322] <= Pix_322[`PIX_WIDTH-1:0];
    Pixels[323] <= Pix_323[`PIX_WIDTH-1:0];
    Pixels[324] <= Pix_324[`PIX_WIDTH-1:0];
    Pixels[325] <= Pix_325[`PIX_WIDTH-1:0];
    Pixels[326] <= Pix_326[`PIX_WIDTH-1:0];
    Pixels[327] <= Pix_327[`PIX_WIDTH-1:0];
    Pixels[328] <= Pix_328[`PIX_WIDTH-1:0];
    Pixels[329] <= Pix_329[`PIX_WIDTH-1:0];
    Pixels[330] <= Pix_330[`PIX_WIDTH-1:0];
    Pixels[331] <= Pix_331[`PIX_WIDTH-1:0];
    Pixels[332] <= Pix_332[`PIX_WIDTH-1:0];
    Pixels[333] <= Pix_333[`PIX_WIDTH-1:0];
    Pixels[334] <= Pix_334[`PIX_WIDTH-1:0];
    Pixels[335] <= Pix_335[`PIX_WIDTH-1:0];
    Pixels[336] <= Pix_336[`PIX_WIDTH-1:0];
    Pixels[337] <= Pix_337[`PIX_WIDTH-1:0];
    Pixels[338] <= Pix_338[`PIX_WIDTH-1:0];
    Pixels[339] <= Pix_339[`PIX_WIDTH-1:0];
    Pixels[340] <= Pix_340[`PIX_WIDTH-1:0];
    Pixels[341] <= Pix_341[`PIX_WIDTH-1:0];
    Pixels[342] <= Pix_342[`PIX_WIDTH-1:0];
    Pixels[343] <= Pix_343[`PIX_WIDTH-1:0];
    Pixels[344] <= Pix_344[`PIX_WIDTH-1:0];
    Pixels[345] <= Pix_345[`PIX_WIDTH-1:0];
    Pixels[346] <= Pix_346[`PIX_WIDTH-1:0];
    Pixels[347] <= Pix_347[`PIX_WIDTH-1:0];
    Pixels[348] <= Pix_348[`PIX_WIDTH-1:0];
    Pixels[349] <= Pix_349[`PIX_WIDTH-1:0];
    Pixels[350] <= Pix_350[`PIX_WIDTH-1:0];
    Pixels[351] <= Pix_351[`PIX_WIDTH-1:0];
    Pixels[352] <= Pix_352[`PIX_WIDTH-1:0];
    Pixels[353] <= Pix_353[`PIX_WIDTH-1:0];
    Pixels[354] <= Pix_354[`PIX_WIDTH-1:0];
    Pixels[355] <= Pix_355[`PIX_WIDTH-1:0];
    Pixels[356] <= Pix_356[`PIX_WIDTH-1:0];
    Pixels[357] <= Pix_357[`PIX_WIDTH-1:0];
    Pixels[358] <= Pix_358[`PIX_WIDTH-1:0];
    Pixels[359] <= Pix_359[`PIX_WIDTH-1:0];
    Pixels[360] <= Pix_360[`PIX_WIDTH-1:0];
    Pixels[361] <= Pix_361[`PIX_WIDTH-1:0];
    Pixels[362] <= Pix_362[`PIX_WIDTH-1:0];
    Pixels[363] <= Pix_363[`PIX_WIDTH-1:0];
    Pixels[364] <= Pix_364[`PIX_WIDTH-1:0];
    Pixels[365] <= Pix_365[`PIX_WIDTH-1:0];
    Pixels[366] <= Pix_366[`PIX_WIDTH-1:0];
    Pixels[367] <= Pix_367[`PIX_WIDTH-1:0];
    Pixels[368] <= Pix_368[`PIX_WIDTH-1:0];
    Pixels[369] <= Pix_369[`PIX_WIDTH-1:0];
    Pixels[370] <= Pix_370[`PIX_WIDTH-1:0];
    Pixels[371] <= Pix_371[`PIX_WIDTH-1:0];
    Pixels[372] <= Pix_372[`PIX_WIDTH-1:0];
    Pixels[373] <= Pix_373[`PIX_WIDTH-1:0];
    Pixels[374] <= Pix_374[`PIX_WIDTH-1:0];
    Pixels[375] <= Pix_375[`PIX_WIDTH-1:0];
    Pixels[376] <= Pix_376[`PIX_WIDTH-1:0];
    Pixels[377] <= Pix_377[`PIX_WIDTH-1:0];
    Pixels[378] <= Pix_378[`PIX_WIDTH-1:0];
    Pixels[379] <= Pix_379[`PIX_WIDTH-1:0];
    Pixels[380] <= Pix_380[`PIX_WIDTH-1:0];
    Pixels[381] <= Pix_381[`PIX_WIDTH-1:0];
    Pixels[382] <= Pix_382[`PIX_WIDTH-1:0];
    Pixels[383] <= Pix_383[`PIX_WIDTH-1:0];
    Pixels[384] <= Pix_384[`PIX_WIDTH-1:0];
    Pixels[385] <= Pix_385[`PIX_WIDTH-1:0];
    Pixels[386] <= Pix_386[`PIX_WIDTH-1:0];
    Pixels[387] <= Pix_387[`PIX_WIDTH-1:0];
    Pixels[388] <= Pix_388[`PIX_WIDTH-1:0];
    Pixels[389] <= Pix_389[`PIX_WIDTH-1:0];
    Pixels[390] <= Pix_390[`PIX_WIDTH-1:0];
    Pixels[391] <= Pix_391[`PIX_WIDTH-1:0];
    Pixels[392] <= Pix_392[`PIX_WIDTH-1:0];
    Pixels[393] <= Pix_393[`PIX_WIDTH-1:0];
    Pixels[394] <= Pix_394[`PIX_WIDTH-1:0];
    Pixels[395] <= Pix_395[`PIX_WIDTH-1:0];
    Pixels[396] <= Pix_396[`PIX_WIDTH-1:0];
    Pixels[397] <= Pix_397[`PIX_WIDTH-1:0];
    Pixels[398] <= Pix_398[`PIX_WIDTH-1:0];
    Pixels[399] <= Pix_399[`PIX_WIDTH-1:0];
    Pixels[400] <= Pix_400[`PIX_WIDTH-1:0];
    Pixels[401] <= Pix_401[`PIX_WIDTH-1:0];
    Pixels[402] <= Pix_402[`PIX_WIDTH-1:0];
    Pixels[403] <= Pix_403[`PIX_WIDTH-1:0];
    Pixels[404] <= Pix_404[`PIX_WIDTH-1:0];
    Pixels[405] <= Pix_405[`PIX_WIDTH-1:0];
    Pixels[406] <= Pix_406[`PIX_WIDTH-1:0];
    Pixels[407] <= Pix_407[`PIX_WIDTH-1:0];
    Pixels[408] <= Pix_408[`PIX_WIDTH-1:0];
    Pixels[409] <= Pix_409[`PIX_WIDTH-1:0];
    Pixels[410] <= Pix_410[`PIX_WIDTH-1:0];
    Pixels[411] <= Pix_411[`PIX_WIDTH-1:0];
    Pixels[412] <= Pix_412[`PIX_WIDTH-1:0];
    Pixels[413] <= Pix_413[`PIX_WIDTH-1:0];
    Pixels[414] <= Pix_414[`PIX_WIDTH-1:0];
    Pixels[415] <= Pix_415[`PIX_WIDTH-1:0];
    Pixels[416] <= Pix_416[`PIX_WIDTH-1:0];
    Pixels[417] <= Pix_417[`PIX_WIDTH-1:0];
    Pixels[418] <= Pix_418[`PIX_WIDTH-1:0];
    Pixels[419] <= Pix_419[`PIX_WIDTH-1:0];
    Pixels[420] <= Pix_420[`PIX_WIDTH-1:0];
    Pixels[421] <= Pix_421[`PIX_WIDTH-1:0];
    Pixels[422] <= Pix_422[`PIX_WIDTH-1:0];
    Pixels[423] <= Pix_423[`PIX_WIDTH-1:0];
    Pixels[424] <= Pix_424[`PIX_WIDTH-1:0];
    Pixels[425] <= Pix_425[`PIX_WIDTH-1:0];
    Pixels[426] <= Pix_426[`PIX_WIDTH-1:0];
    Pixels[427] <= Pix_427[`PIX_WIDTH-1:0];
    Pixels[428] <= Pix_428[`PIX_WIDTH-1:0];
    Pixels[429] <= Pix_429[`PIX_WIDTH-1:0];
    Pixels[430] <= Pix_430[`PIX_WIDTH-1:0];
    Pixels[431] <= Pix_431[`PIX_WIDTH-1:0];
    Pixels[432] <= Pix_432[`PIX_WIDTH-1:0];
    Pixels[433] <= Pix_433[`PIX_WIDTH-1:0];
    Pixels[434] <= Pix_434[`PIX_WIDTH-1:0];
    Pixels[435] <= Pix_435[`PIX_WIDTH-1:0];
    Pixels[436] <= Pix_436[`PIX_WIDTH-1:0];
    Pixels[437] <= Pix_437[`PIX_WIDTH-1:0];
    Pixels[438] <= Pix_438[`PIX_WIDTH-1:0];
    Pixels[439] <= Pix_439[`PIX_WIDTH-1:0];
    Pixels[440] <= Pix_440[`PIX_WIDTH-1:0];
    Pixels[441] <= Pix_441[`PIX_WIDTH-1:0];
    Pixels[442] <= Pix_442[`PIX_WIDTH-1:0];
    Pixels[443] <= Pix_443[`PIX_WIDTH-1:0];
    Pixels[444] <= Pix_444[`PIX_WIDTH-1:0];
    Pixels[445] <= Pix_445[`PIX_WIDTH-1:0];
    Pixels[446] <= Pix_446[`PIX_WIDTH-1:0];
    Pixels[447] <= Pix_447[`PIX_WIDTH-1:0];
    Pixels[448] <= Pix_448[`PIX_WIDTH-1:0];
    Pixels[449] <= Pix_449[`PIX_WIDTH-1:0];
    Pixels[450] <= Pix_450[`PIX_WIDTH-1:0];
    Pixels[451] <= Pix_451[`PIX_WIDTH-1:0];
    Pixels[452] <= Pix_452[`PIX_WIDTH-1:0];
    Pixels[453] <= Pix_453[`PIX_WIDTH-1:0];
    Pixels[454] <= Pix_454[`PIX_WIDTH-1:0];
    Pixels[455] <= Pix_455[`PIX_WIDTH-1:0];
    Pixels[456] <= Pix_456[`PIX_WIDTH-1:0];
    Pixels[457] <= Pix_457[`PIX_WIDTH-1:0];
    Pixels[458] <= Pix_458[`PIX_WIDTH-1:0];
    Pixels[459] <= Pix_459[`PIX_WIDTH-1:0];
    Pixels[460] <= Pix_460[`PIX_WIDTH-1:0];
    Pixels[461] <= Pix_461[`PIX_WIDTH-1:0];
    Pixels[462] <= Pix_462[`PIX_WIDTH-1:0];
    Pixels[463] <= Pix_463[`PIX_WIDTH-1:0];
    Pixels[464] <= Pix_464[`PIX_WIDTH-1:0];
    Pixels[465] <= Pix_465[`PIX_WIDTH-1:0];
    Pixels[466] <= Pix_466[`PIX_WIDTH-1:0];
    Pixels[467] <= Pix_467[`PIX_WIDTH-1:0];
    Pixels[468] <= Pix_468[`PIX_WIDTH-1:0];
    Pixels[469] <= Pix_469[`PIX_WIDTH-1:0];
    Pixels[470] <= Pix_470[`PIX_WIDTH-1:0];
    Pixels[471] <= Pix_471[`PIX_WIDTH-1:0];
    Pixels[472] <= Pix_472[`PIX_WIDTH-1:0];
    Pixels[473] <= Pix_473[`PIX_WIDTH-1:0];
    Pixels[474] <= Pix_474[`PIX_WIDTH-1:0];
    Pixels[475] <= Pix_475[`PIX_WIDTH-1:0];
    Pixels[476] <= Pix_476[`PIX_WIDTH-1:0];
    Pixels[477] <= Pix_477[`PIX_WIDTH-1:0];
    Pixels[478] <= Pix_478[`PIX_WIDTH-1:0];
    Pixels[479] <= Pix_479[`PIX_WIDTH-1:0];
    Pixels[480] <= Pix_480[`PIX_WIDTH-1:0];
    Pixels[481] <= Pix_481[`PIX_WIDTH-1:0];
    Pixels[482] <= Pix_482[`PIX_WIDTH-1:0];
    Pixels[483] <= Pix_483[`PIX_WIDTH-1:0];
    Pixels[484] <= Pix_484[`PIX_WIDTH-1:0];
    Pixels[485] <= Pix_485[`PIX_WIDTH-1:0];
    Pixels[486] <= Pix_486[`PIX_WIDTH-1:0];
    Pixels[487] <= Pix_487[`PIX_WIDTH-1:0];
    Pixels[488] <= Pix_488[`PIX_WIDTH-1:0];
    Pixels[489] <= Pix_489[`PIX_WIDTH-1:0];
    Pixels[490] <= Pix_490[`PIX_WIDTH-1:0];
    Pixels[491] <= Pix_491[`PIX_WIDTH-1:0];
    Pixels[492] <= Pix_492[`PIX_WIDTH-1:0];
    Pixels[493] <= Pix_493[`PIX_WIDTH-1:0];
    Pixels[494] <= Pix_494[`PIX_WIDTH-1:0];
    Pixels[495] <= Pix_495[`PIX_WIDTH-1:0];
    Pixels[496] <= Pix_496[`PIX_WIDTH-1:0];
    Pixels[497] <= Pix_497[`PIX_WIDTH-1:0];
    Pixels[498] <= Pix_498[`PIX_WIDTH-1:0];
    Pixels[499] <= Pix_499[`PIX_WIDTH-1:0];
    Pixels[500] <= Pix_500[`PIX_WIDTH-1:0];
    Pixels[501] <= Pix_501[`PIX_WIDTH-1:0];
    Pixels[502] <= Pix_502[`PIX_WIDTH-1:0];
    Pixels[503] <= Pix_503[`PIX_WIDTH-1:0];
    Pixels[504] <= Pix_504[`PIX_WIDTH-1:0];
    Pixels[505] <= Pix_505[`PIX_WIDTH-1:0];
    Pixels[506] <= Pix_506[`PIX_WIDTH-1:0];
    Pixels[507] <= Pix_507[`PIX_WIDTH-1:0];
    Pixels[508] <= Pix_508[`PIX_WIDTH-1:0];
    Pixels[509] <= Pix_509[`PIX_WIDTH-1:0];
    Pixels[510] <= Pix_510[`PIX_WIDTH-1:0];
    Pixels[511] <= Pix_511[`PIX_WIDTH-1:0];
    Pixels[512] <= Pix_512[`PIX_WIDTH-1:0];
    Pixels[513] <= Pix_513[`PIX_WIDTH-1:0];
    Pixels[514] <= Pix_514[`PIX_WIDTH-1:0];
    Pixels[515] <= Pix_515[`PIX_WIDTH-1:0];
    Pixels[516] <= Pix_516[`PIX_WIDTH-1:0];
    Pixels[517] <= Pix_517[`PIX_WIDTH-1:0];
    Pixels[518] <= Pix_518[`PIX_WIDTH-1:0];
    Pixels[519] <= Pix_519[`PIX_WIDTH-1:0];
    Pixels[520] <= Pix_520[`PIX_WIDTH-1:0];
    Pixels[521] <= Pix_521[`PIX_WIDTH-1:0];
    Pixels[522] <= Pix_522[`PIX_WIDTH-1:0];
    Pixels[523] <= Pix_523[`PIX_WIDTH-1:0];
    Pixels[524] <= Pix_524[`PIX_WIDTH-1:0];
    Pixels[525] <= Pix_525[`PIX_WIDTH-1:0];
    Pixels[526] <= Pix_526[`PIX_WIDTH-1:0];
    Pixels[527] <= Pix_527[`PIX_WIDTH-1:0];
    Pixels[528] <= Pix_528[`PIX_WIDTH-1:0];
    Pixels[529] <= Pix_529[`PIX_WIDTH-1:0];
    Pixels[530] <= Pix_530[`PIX_WIDTH-1:0];
    Pixels[531] <= Pix_531[`PIX_WIDTH-1:0];
    Pixels[532] <= Pix_532[`PIX_WIDTH-1:0];
    Pixels[533] <= Pix_533[`PIX_WIDTH-1:0];
    Pixels[534] <= Pix_534[`PIX_WIDTH-1:0];
    Pixels[535] <= Pix_535[`PIX_WIDTH-1:0];
    Pixels[536] <= Pix_536[`PIX_WIDTH-1:0];
    Pixels[537] <= Pix_537[`PIX_WIDTH-1:0];
    Pixels[538] <= Pix_538[`PIX_WIDTH-1:0];
    Pixels[539] <= Pix_539[`PIX_WIDTH-1:0];
    Pixels[540] <= Pix_540[`PIX_WIDTH-1:0];
    Pixels[541] <= Pix_541[`PIX_WIDTH-1:0];
    Pixels[542] <= Pix_542[`PIX_WIDTH-1:0];
    Pixels[543] <= Pix_543[`PIX_WIDTH-1:0];
    Pixels[544] <= Pix_544[`PIX_WIDTH-1:0];
    Pixels[545] <= Pix_545[`PIX_WIDTH-1:0];
    Pixels[546] <= Pix_546[`PIX_WIDTH-1:0];
    Pixels[547] <= Pix_547[`PIX_WIDTH-1:0];
    Pixels[548] <= Pix_548[`PIX_WIDTH-1:0];
    Pixels[549] <= Pix_549[`PIX_WIDTH-1:0];
    Pixels[550] <= Pix_550[`PIX_WIDTH-1:0];
    Pixels[551] <= Pix_551[`PIX_WIDTH-1:0];
    Pixels[552] <= Pix_552[`PIX_WIDTH-1:0];
    Pixels[553] <= Pix_553[`PIX_WIDTH-1:0];
    Pixels[554] <= Pix_554[`PIX_WIDTH-1:0];
    Pixels[555] <= Pix_555[`PIX_WIDTH-1:0];
    Pixels[556] <= Pix_556[`PIX_WIDTH-1:0];
    Pixels[557] <= Pix_557[`PIX_WIDTH-1:0];
    Pixels[558] <= Pix_558[`PIX_WIDTH-1:0];
    Pixels[559] <= Pix_559[`PIX_WIDTH-1:0];
    Pixels[560] <= Pix_560[`PIX_WIDTH-1:0];
    Pixels[561] <= Pix_561[`PIX_WIDTH-1:0];
    Pixels[562] <= Pix_562[`PIX_WIDTH-1:0];
    Pixels[563] <= Pix_563[`PIX_WIDTH-1:0];
    Pixels[564] <= Pix_564[`PIX_WIDTH-1:0];
    Pixels[565] <= Pix_565[`PIX_WIDTH-1:0];
    Pixels[566] <= Pix_566[`PIX_WIDTH-1:0];
    Pixels[567] <= Pix_567[`PIX_WIDTH-1:0];
    Pixels[568] <= Pix_568[`PIX_WIDTH-1:0];
    Pixels[569] <= Pix_569[`PIX_WIDTH-1:0];
    Pixels[570] <= Pix_570[`PIX_WIDTH-1:0];
    Pixels[571] <= Pix_571[`PIX_WIDTH-1:0];
    Pixels[572] <= Pix_572[`PIX_WIDTH-1:0];
    Pixels[573] <= Pix_573[`PIX_WIDTH-1:0];
    Pixels[574] <= Pix_574[`PIX_WIDTH-1:0];
    Pixels[575] <= Pix_575[`PIX_WIDTH-1:0];
    Pixels[576] <= Pix_576[`PIX_WIDTH-1:0];
    Pixels[577] <= Pix_577[`PIX_WIDTH-1:0];
    Pixels[578] <= Pix_578[`PIX_WIDTH-1:0];
    Pixels[579] <= Pix_579[`PIX_WIDTH-1:0];
    Pixels[580] <= Pix_580[`PIX_WIDTH-1:0];
    Pixels[581] <= Pix_581[`PIX_WIDTH-1:0];
    Pixels[582] <= Pix_582[`PIX_WIDTH-1:0];
    Pixels[583] <= Pix_583[`PIX_WIDTH-1:0];
    Pixels[584] <= Pix_584[`PIX_WIDTH-1:0];
    Pixels[585] <= Pix_585[`PIX_WIDTH-1:0];
    Pixels[586] <= Pix_586[`PIX_WIDTH-1:0];
    Pixels[587] <= Pix_587[`PIX_WIDTH-1:0];
    Pixels[588] <= Pix_588[`PIX_WIDTH-1:0];
    Pixels[589] <= Pix_589[`PIX_WIDTH-1:0];
    Pixels[590] <= Pix_590[`PIX_WIDTH-1:0];
    Pixels[591] <= Pix_591[`PIX_WIDTH-1:0];
    Pixels[592] <= Pix_592[`PIX_WIDTH-1:0];
    Pixels[593] <= Pix_593[`PIX_WIDTH-1:0];
    Pixels[594] <= Pix_594[`PIX_WIDTH-1:0];
    Pixels[595] <= Pix_595[`PIX_WIDTH-1:0];
    Pixels[596] <= Pix_596[`PIX_WIDTH-1:0];
    Pixels[597] <= Pix_597[`PIX_WIDTH-1:0];
    Pixels[598] <= Pix_598[`PIX_WIDTH-1:0];
    Pixels[599] <= Pix_599[`PIX_WIDTH-1:0];
    Pixels[600] <= Pix_600[`PIX_WIDTH-1:0];
    Pixels[601] <= Pix_601[`PIX_WIDTH-1:0];
    Pixels[602] <= Pix_602[`PIX_WIDTH-1:0];
    Pixels[603] <= Pix_603[`PIX_WIDTH-1:0];
    Pixels[604] <= Pix_604[`PIX_WIDTH-1:0];
    Pixels[605] <= Pix_605[`PIX_WIDTH-1:0];
    Pixels[606] <= Pix_606[`PIX_WIDTH-1:0];
    Pixels[607] <= Pix_607[`PIX_WIDTH-1:0];
    Pixels[608] <= Pix_608[`PIX_WIDTH-1:0];
    Pixels[609] <= Pix_609[`PIX_WIDTH-1:0];
    Pixels[610] <= Pix_610[`PIX_WIDTH-1:0];
    Pixels[611] <= Pix_611[`PIX_WIDTH-1:0];
    Pixels[612] <= Pix_612[`PIX_WIDTH-1:0];
    Pixels[613] <= Pix_613[`PIX_WIDTH-1:0];
    Pixels[614] <= Pix_614[`PIX_WIDTH-1:0];
    Pixels[615] <= Pix_615[`PIX_WIDTH-1:0];
    Pixels[616] <= Pix_616[`PIX_WIDTH-1:0];
    Pixels[617] <= Pix_617[`PIX_WIDTH-1:0];
    Pixels[618] <= Pix_618[`PIX_WIDTH-1:0];
    Pixels[619] <= Pix_619[`PIX_WIDTH-1:0];
    Pixels[620] <= Pix_620[`PIX_WIDTH-1:0];
    Pixels[621] <= Pix_621[`PIX_WIDTH-1:0];
    Pixels[622] <= Pix_622[`PIX_WIDTH-1:0];
    Pixels[623] <= Pix_623[`PIX_WIDTH-1:0];
    Pixels[624] <= Pix_624[`PIX_WIDTH-1:0];
    Pixels[625] <= Pix_625[`PIX_WIDTH-1:0];
    Pixels[626] <= Pix_626[`PIX_WIDTH-1:0];
    Pixels[627] <= Pix_627[`PIX_WIDTH-1:0];
    Pixels[628] <= Pix_628[`PIX_WIDTH-1:0];
    Pixels[629] <= Pix_629[`PIX_WIDTH-1:0];
    Pixels[630] <= Pix_630[`PIX_WIDTH-1:0];
    Pixels[631] <= Pix_631[`PIX_WIDTH-1:0];
    Pixels[632] <= Pix_632[`PIX_WIDTH-1:0];
    Pixels[633] <= Pix_633[`PIX_WIDTH-1:0];
    Pixels[634] <= Pix_634[`PIX_WIDTH-1:0];
    Pixels[635] <= Pix_635[`PIX_WIDTH-1:0];
    Pixels[636] <= Pix_636[`PIX_WIDTH-1:0];
    Pixels[637] <= Pix_637[`PIX_WIDTH-1:0];
    Pixels[638] <= Pix_638[`PIX_WIDTH-1:0];
    Pixels[639] <= Pix_639[`PIX_WIDTH-1:0];
    Pixels[640] <= Pix_640[`PIX_WIDTH-1:0];
    Pixels[641] <= Pix_641[`PIX_WIDTH-1:0];
    Pixels[642] <= Pix_642[`PIX_WIDTH-1:0];
    Pixels[643] <= Pix_643[`PIX_WIDTH-1:0];
    Pixels[644] <= Pix_644[`PIX_WIDTH-1:0];
    Pixels[645] <= Pix_645[`PIX_WIDTH-1:0];
    Pixels[646] <= Pix_646[`PIX_WIDTH-1:0];
    Pixels[647] <= Pix_647[`PIX_WIDTH-1:0];
    Pixels[648] <= Pix_648[`PIX_WIDTH-1:0];
    Pixels[649] <= Pix_649[`PIX_WIDTH-1:0];
    Pixels[650] <= Pix_650[`PIX_WIDTH-1:0];
    Pixels[651] <= Pix_651[`PIX_WIDTH-1:0];
    Pixels[652] <= Pix_652[`PIX_WIDTH-1:0];
    Pixels[653] <= Pix_653[`PIX_WIDTH-1:0];
    Pixels[654] <= Pix_654[`PIX_WIDTH-1:0];
    Pixels[655] <= Pix_655[`PIX_WIDTH-1:0];
    Pixels[656] <= Pix_656[`PIX_WIDTH-1:0];
    Pixels[657] <= Pix_657[`PIX_WIDTH-1:0];
    Pixels[658] <= Pix_658[`PIX_WIDTH-1:0];
    Pixels[659] <= Pix_659[`PIX_WIDTH-1:0];
    Pixels[660] <= Pix_660[`PIX_WIDTH-1:0];
    Pixels[661] <= Pix_661[`PIX_WIDTH-1:0];
    Pixels[662] <= Pix_662[`PIX_WIDTH-1:0];
    Pixels[663] <= Pix_663[`PIX_WIDTH-1:0];
    Pixels[664] <= Pix_664[`PIX_WIDTH-1:0];
    Pixels[665] <= Pix_665[`PIX_WIDTH-1:0];
    Pixels[666] <= Pix_666[`PIX_WIDTH-1:0];
    Pixels[667] <= Pix_667[`PIX_WIDTH-1:0];
    Pixels[668] <= Pix_668[`PIX_WIDTH-1:0];
    Pixels[669] <= Pix_669[`PIX_WIDTH-1:0];
    Pixels[670] <= Pix_670[`PIX_WIDTH-1:0];
    Pixels[671] <= Pix_671[`PIX_WIDTH-1:0];
    Pixels[672] <= Pix_672[`PIX_WIDTH-1:0];
    Pixels[673] <= Pix_673[`PIX_WIDTH-1:0];
    Pixels[674] <= Pix_674[`PIX_WIDTH-1:0];
    Pixels[675] <= Pix_675[`PIX_WIDTH-1:0];
    Pixels[676] <= Pix_676[`PIX_WIDTH-1:0];
    Pixels[677] <= Pix_677[`PIX_WIDTH-1:0];
    Pixels[678] <= Pix_678[`PIX_WIDTH-1:0];
    Pixels[679] <= Pix_679[`PIX_WIDTH-1:0];
    Pixels[680] <= Pix_680[`PIX_WIDTH-1:0];
    Pixels[681] <= Pix_681[`PIX_WIDTH-1:0];
    Pixels[682] <= Pix_682[`PIX_WIDTH-1:0];
    Pixels[683] <= Pix_683[`PIX_WIDTH-1:0];
    Pixels[684] <= Pix_684[`PIX_WIDTH-1:0];
    Pixels[685] <= Pix_685[`PIX_WIDTH-1:0];
    Pixels[686] <= Pix_686[`PIX_WIDTH-1:0];
    Pixels[687] <= Pix_687[`PIX_WIDTH-1:0];
    Pixels[688] <= Pix_688[`PIX_WIDTH-1:0];
    Pixels[689] <= Pix_689[`PIX_WIDTH-1:0];
    Pixels[690] <= Pix_690[`PIX_WIDTH-1:0];
    Pixels[691] <= Pix_691[`PIX_WIDTH-1:0];
    Pixels[692] <= Pix_692[`PIX_WIDTH-1:0];
    Pixels[693] <= Pix_693[`PIX_WIDTH-1:0];
    Pixels[694] <= Pix_694[`PIX_WIDTH-1:0];
    Pixels[695] <= Pix_695[`PIX_WIDTH-1:0];
    Pixels[696] <= Pix_696[`PIX_WIDTH-1:0];
    Pixels[697] <= Pix_697[`PIX_WIDTH-1:0];
    Pixels[698] <= Pix_698[`PIX_WIDTH-1:0];
    Pixels[699] <= Pix_699[`PIX_WIDTH-1:0];
    Pixels[700] <= Pix_700[`PIX_WIDTH-1:0];
    Pixels[701] <= Pix_701[`PIX_WIDTH-1:0];
    Pixels[702] <= Pix_702[`PIX_WIDTH-1:0];
    Pixels[703] <= Pix_703[`PIX_WIDTH-1:0];
    Pixels[704] <= Pix_704[`PIX_WIDTH-1:0];
    Pixels[705] <= Pix_705[`PIX_WIDTH-1:0];
    Pixels[706] <= Pix_706[`PIX_WIDTH-1:0];
    Pixels[707] <= Pix_707[`PIX_WIDTH-1:0];
    Pixels[708] <= Pix_708[`PIX_WIDTH-1:0];
    Pixels[709] <= Pix_709[`PIX_WIDTH-1:0];
    Pixels[710] <= Pix_710[`PIX_WIDTH-1:0];
    Pixels[711] <= Pix_711[`PIX_WIDTH-1:0];
    Pixels[712] <= Pix_712[`PIX_WIDTH-1:0];
    Pixels[713] <= Pix_713[`PIX_WIDTH-1:0];
    Pixels[714] <= Pix_714[`PIX_WIDTH-1:0];
    Pixels[715] <= Pix_715[`PIX_WIDTH-1:0];
    Pixels[716] <= Pix_716[`PIX_WIDTH-1:0];
    Pixels[717] <= Pix_717[`PIX_WIDTH-1:0];
    Pixels[718] <= Pix_718[`PIX_WIDTH-1:0];
    Pixels[719] <= Pix_719[`PIX_WIDTH-1:0];
    Pixels[720] <= Pix_720[`PIX_WIDTH-1:0];
    Pixels[721] <= Pix_721[`PIX_WIDTH-1:0];
    Pixels[722] <= Pix_722[`PIX_WIDTH-1:0];
    Pixels[723] <= Pix_723[`PIX_WIDTH-1:0];
    Pixels[724] <= Pix_724[`PIX_WIDTH-1:0];
    Pixels[725] <= Pix_725[`PIX_WIDTH-1:0];
    Pixels[726] <= Pix_726[`PIX_WIDTH-1:0];
    Pixels[727] <= Pix_727[`PIX_WIDTH-1:0];
    Pixels[728] <= Pix_728[`PIX_WIDTH-1:0];
    Pixels[729] <= Pix_729[`PIX_WIDTH-1:0];
    Pixels[730] <= Pix_730[`PIX_WIDTH-1:0];
    Pixels[731] <= Pix_731[`PIX_WIDTH-1:0];
    Pixels[732] <= Pix_732[`PIX_WIDTH-1:0];
    Pixels[733] <= Pix_733[`PIX_WIDTH-1:0];
    Pixels[734] <= Pix_734[`PIX_WIDTH-1:0];
    Pixels[735] <= Pix_735[`PIX_WIDTH-1:0];
    Pixels[736] <= Pix_736[`PIX_WIDTH-1:0];
    Pixels[737] <= Pix_737[`PIX_WIDTH-1:0];
    Pixels[738] <= Pix_738[`PIX_WIDTH-1:0];
    Pixels[739] <= Pix_739[`PIX_WIDTH-1:0];
    Pixels[740] <= Pix_740[`PIX_WIDTH-1:0];
    Pixels[741] <= Pix_741[`PIX_WIDTH-1:0];
    Pixels[742] <= Pix_742[`PIX_WIDTH-1:0];
    Pixels[743] <= Pix_743[`PIX_WIDTH-1:0];
    Pixels[744] <= Pix_744[`PIX_WIDTH-1:0];
    Pixels[745] <= Pix_745[`PIX_WIDTH-1:0];
    Pixels[746] <= Pix_746[`PIX_WIDTH-1:0];
    Pixels[747] <= Pix_747[`PIX_WIDTH-1:0];
    Pixels[748] <= Pix_748[`PIX_WIDTH-1:0];
    Pixels[749] <= Pix_749[`PIX_WIDTH-1:0];
    Pixels[750] <= Pix_750[`PIX_WIDTH-1:0];
    Pixels[751] <= Pix_751[`PIX_WIDTH-1:0];
    Pixels[752] <= Pix_752[`PIX_WIDTH-1:0];
    Pixels[753] <= Pix_753[`PIX_WIDTH-1:0];
    Pixels[754] <= Pix_754[`PIX_WIDTH-1:0];
    Pixels[755] <= Pix_755[`PIX_WIDTH-1:0];
    Pixels[756] <= Pix_756[`PIX_WIDTH-1:0];
    Pixels[757] <= Pix_757[`PIX_WIDTH-1:0];
    Pixels[758] <= Pix_758[`PIX_WIDTH-1:0];
    Pixels[759] <= Pix_759[`PIX_WIDTH-1:0];
    Pixels[760] <= Pix_760[`PIX_WIDTH-1:0];
    Pixels[761] <= Pix_761[`PIX_WIDTH-1:0];
    Pixels[762] <= Pix_762[`PIX_WIDTH-1:0];
    Pixels[763] <= Pix_763[`PIX_WIDTH-1:0];
    Pixels[764] <= Pix_764[`PIX_WIDTH-1:0];
    Pixels[765] <= Pix_765[`PIX_WIDTH-1:0];
    Pixels[766] <= Pix_766[`PIX_WIDTH-1:0];
    Pixels[767] <= Pix_767[`PIX_WIDTH-1:0];
    Pixels[768] <= Pix_768[`PIX_WIDTH-1:0];
    Pixels[769] <= Pix_769[`PIX_WIDTH-1:0];
    Pixels[770] <= Pix_770[`PIX_WIDTH-1:0];
    Pixels[771] <= Pix_771[`PIX_WIDTH-1:0];
    Pixels[772] <= Pix_772[`PIX_WIDTH-1:0];
    Pixels[773] <= Pix_773[`PIX_WIDTH-1:0];
    Pixels[774] <= Pix_774[`PIX_WIDTH-1:0];
    Pixels[775] <= Pix_775[`PIX_WIDTH-1:0];
    Pixels[776] <= Pix_776[`PIX_WIDTH-1:0];
    Pixels[777] <= Pix_777[`PIX_WIDTH-1:0];
    Pixels[778] <= Pix_778[`PIX_WIDTH-1:0];
    Pixels[779] <= Pix_779[`PIX_WIDTH-1:0];
    Pixels[780] <= Pix_780[`PIX_WIDTH-1:0];
    Pixels[781] <= Pix_781[`PIX_WIDTH-1:0];
    Pixels[782] <= Pix_782[`PIX_WIDTH-1:0];
    Pixels[783] <= Pix_783[`PIX_WIDTH-1:0];
    Pixels[784] <= Pix_784[`PIX_WIDTH-1:0]; // always 1, Weights[784] = bias
end

// internal regs
reg neuron_en_r; // neuron enable 
reg neuron_reset_r; // neuron reset
reg max_en_r; // enable max selector
reg max_reset_r; // max selector reset
// reg [`PIX_WIDTH-1:0] count_r; // counter

reg [5:0] select_count;

// neuron_0 
wire [`PIX_WIDTH-1:0] pixel0_0,pixel0_1,pixel0_2,pixel0_3,pixel0_4,pixel0_5,pixel0_6,pixel0_7,pixel0_8,pixel0_9,pixel0_10,pixel0_11,pixel0_12,pixel0_13,pixel0_14,pixel0_15;
Pixel_MUX pixel_mux0_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel0_0));
Pixel_MUX pixel_mux0_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_1));
Pixel_MUX pixel_mux0_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_2));
Pixel_MUX pixel_mux0_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_3));
Pixel_MUX pixel_mux0_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_4));
Pixel_MUX pixel_mux0_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_5));
Pixel_MUX pixel_mux0_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_6));
Pixel_MUX pixel_mux0_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_7));
Pixel_MUX pixel_mux0_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_8));
Pixel_MUX pixel_mux0_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_9));
Pixel_MUX pixel_mux0_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_10));
Pixel_MUX pixel_mux0_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_11));
Pixel_MUX pixel_mux0_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_12));
Pixel_MUX pixel_mux0_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_13));
Pixel_MUX pixel_mux0_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_14));
Pixel_MUX pixel_mux0_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel0_15));
wire [`WGT_WIDTH-1:0] weight0_0,weight0_1,weight0_2,weight0_3,weight0_4,weight0_5,weight0_6,weight0_7,weight0_8,weight0_9,weight0_10,weight0_11,weight0_12,weight0_13,weight0_14,weight0_15;
Weight_MUX weight_mux0_0(.Weight_0(Wgt_0_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_0_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight0_0));
Weight_MUX weight_mux0_1(.Weight_0(Wgt_0_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_1));
Weight_MUX weight_mux0_2(.Weight_0(Wgt_0_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_2));
Weight_MUX weight_mux0_3(.Weight_0(Wgt_0_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_3));
Weight_MUX weight_mux0_4(.Weight_0(Wgt_0_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_4));
Weight_MUX weight_mux0_5(.Weight_0(Wgt_0_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_5));
Weight_MUX weight_mux0_6(.Weight_0(Wgt_0_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_6));
Weight_MUX weight_mux0_7(.Weight_0(Wgt_0_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_7));
Weight_MUX weight_mux0_8(.Weight_0(Wgt_0_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_8));
Weight_MUX weight_mux0_9(.Weight_0(Wgt_0_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_9));
Weight_MUX weight_mux0_10(.Weight_0(Wgt_0_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_10));
Weight_MUX weight_mux0_11(.Weight_0(Wgt_0_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_11));
Weight_MUX weight_mux0_12(.Weight_0(Wgt_0_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_12));
Weight_MUX weight_mux0_13(.Weight_0(Wgt_0_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_13));
Weight_MUX weight_mux0_14(.Weight_0(Wgt_0_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_14));
Weight_MUX weight_mux0_15(.Weight_0(Wgt_0_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_0_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_0_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_0_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_0_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_0_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_0_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_0_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_0_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_0_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_0_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_0_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_0_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_0_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_0_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_0_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_0_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_0_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_0_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_0_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_0_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_0_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_0_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_0_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_0_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_0_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_0_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_0_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_0_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_0_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_0_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_0_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_0_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_0_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_0_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_0_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_0_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_0_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_0_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_0_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_0_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_0_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_0_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_0_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_0_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_0_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_0_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_0_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_0_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight0_15));
wire [25:0] out_n0;
Neuron neuron_0(.Weight_0(weight0_0),.Weight_1(weight0_1),.Weight_2(weight0_2),.Weight_3(weight0_3),.Weight_4(weight0_4),.Weight_5(weight0_5),.Weight_6(weight0_6),.Weight_7(weight0_7),.Weight_8(weight0_8),.Weight_9(weight0_9),.Weight_10(weight0_10),.Weight_11(weight0_11),.Weight_12(weight0_12),.Weight_13(weight0_13),.Weight_14(weight0_14),.Weight_15(weight0_15),.Pixel_0(pixel0_0),.Pixel_1(pixel0_1),.Pixel_2(pixel0_2),.Pixel_3(pixel0_3),.Pixel_4(pixel0_4),.Pixel_5(pixel0_5),.Pixel_6(pixel0_6),.Pixel_7(pixel0_7),.Pixel_8(pixel0_8),.Pixel_9(pixel0_9),.Pixel_10(pixel0_10),.Pixel_11(pixel0_11),.Pixel_12(pixel0_12),.Pixel_13(pixel0_13),.Pixel_14(pixel0_14),.Pixel_15(pixel0_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n0));

// neuron_1
wire [`PIX_WIDTH-1:0] pixel1_0,pixel1_1,pixel1_2,pixel1_3,pixel1_4,pixel1_5,pixel1_6,pixel1_7,pixel1_8,pixel1_9,pixel1_10,pixel1_11,pixel1_12,pixel1_13,pixel1_14,pixel1_15;
Pixel_MUX pixel_mux1_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel1_0));
Pixel_MUX pixel_mux1_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_1));
Pixel_MUX pixel_mux1_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_2));
Pixel_MUX pixel_mux1_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_3));
Pixel_MUX pixel_mux1_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_4));
Pixel_MUX pixel_mux1_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_5));
Pixel_MUX pixel_mux1_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_6));
Pixel_MUX pixel_mux1_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_7));
Pixel_MUX pixel_mux1_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_8));
Pixel_MUX pixel_mux1_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_9));
Pixel_MUX pixel_mux1_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_10));
Pixel_MUX pixel_mux1_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_11));
Pixel_MUX pixel_mux1_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_12));
Pixel_MUX pixel_mux1_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_13));
Pixel_MUX pixel_mux1_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_14));
Pixel_MUX pixel_mux1_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel1_15));
wire [`WGT_WIDTH-1:0] weight1_0,weight1_1,weight1_2,weight1_3,weight1_4,weight1_5,weight1_6,weight1_7,weight1_8,weight1_9,weight1_10,weight1_11,weight1_12,weight1_13,weight1_14,weight1_15;
Weight_MUX weight_mux1_0(.Weight_0(Wgt_1_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_1_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight1_0));
Weight_MUX weight_mux1_1(.Weight_0(Wgt_1_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_1));
Weight_MUX weight_mux1_2(.Weight_0(Wgt_1_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_2));
Weight_MUX weight_mux1_3(.Weight_0(Wgt_1_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_3));
Weight_MUX weight_mux1_4(.Weight_0(Wgt_1_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_4));
Weight_MUX weight_mux1_5(.Weight_0(Wgt_1_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_5));
Weight_MUX weight_mux1_6(.Weight_0(Wgt_1_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_6));
Weight_MUX weight_mux1_7(.Weight_0(Wgt_1_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_7));
Weight_MUX weight_mux1_8(.Weight_0(Wgt_1_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_8));
Weight_MUX weight_mux1_9(.Weight_0(Wgt_1_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_9));
Weight_MUX weight_mux1_10(.Weight_0(Wgt_1_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_10));
Weight_MUX weight_mux1_11(.Weight_0(Wgt_1_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_11));
Weight_MUX weight_mux1_12(.Weight_0(Wgt_1_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_12));
Weight_MUX weight_mux1_13(.Weight_0(Wgt_1_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_13));
Weight_MUX weight_mux1_14(.Weight_0(Wgt_1_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_14));
Weight_MUX weight_mux1_15(.Weight_0(Wgt_1_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_1_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_1_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_1_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_1_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_1_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_1_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_1_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_1_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_1_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_1_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_1_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_1_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_1_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_1_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_1_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_1_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_1_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_1_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_1_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_1_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_1_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_1_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_1_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_1_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_1_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_1_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_1_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_1_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_1_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_1_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_1_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_1_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_1_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_1_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_1_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_1_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_1_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_1_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_1_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_1_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_1_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_1_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_1_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_1_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_1_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_1_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_1_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_1_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight1_15));
wire [25:0] out_n1;
Neuron neuron_1(.Weight_0(weight1_0),.Weight_1(weight1_1),.Weight_2(weight1_2),.Weight_3(weight1_3),.Weight_4(weight1_4),.Weight_5(weight1_5),.Weight_6(weight1_6),.Weight_7(weight1_7),.Weight_8(weight1_8),.Weight_9(weight1_9),.Weight_10(weight1_10),.Weight_11(weight1_11),.Weight_12(weight1_12),.Weight_13(weight1_13),.Weight_14(weight1_14),.Weight_15(weight1_15),.Pixel_0(pixel1_0),.Pixel_1(pixel1_1),.Pixel_2(pixel1_2),.Pixel_3(pixel1_3),.Pixel_4(pixel1_4),.Pixel_5(pixel1_5),.Pixel_6(pixel1_6),.Pixel_7(pixel1_7),.Pixel_8(pixel1_8),.Pixel_9(pixel1_9),.Pixel_10(pixel1_10),.Pixel_11(pixel1_11),.Pixel_12(pixel1_12),.Pixel_13(pixel1_13),.Pixel_14(pixel1_14),.Pixel_15(pixel1_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n1));

// neuron_2
wire [`PIX_WIDTH-1:0] pixel2_0,pixel2_1,pixel2_2,pixel2_3,pixel2_4,pixel2_5,pixel2_6,pixel2_7,pixel2_8,pixel2_9,pixel2_10,pixel2_11,pixel2_12,pixel2_13,pixel2_14,pixel2_15;
Pixel_MUX pixel_mux2_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel2_0));
Pixel_MUX pixel_mux2_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_1));
Pixel_MUX pixel_mux2_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_2));
Pixel_MUX pixel_mux2_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_3));
Pixel_MUX pixel_mux2_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_4));
Pixel_MUX pixel_mux2_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_5));
Pixel_MUX pixel_mux2_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_6));
Pixel_MUX pixel_mux2_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_7));
Pixel_MUX pixel_mux2_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_8));
Pixel_MUX pixel_mux2_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_9));
Pixel_MUX pixel_mux2_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_10));
Pixel_MUX pixel_mux2_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_11));
Pixel_MUX pixel_mux2_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_12));
Pixel_MUX pixel_mux2_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_13));
Pixel_MUX pixel_mux2_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_14));
Pixel_MUX pixel_mux2_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel2_15));
wire [`WGT_WIDTH-1:0] weight2_0,weight2_1,weight2_2,weight2_3,weight2_4,weight2_5,weight2_6,weight2_7,weight2_8,weight2_9,weight2_10,weight2_11,weight2_12,weight2_13,weight2_14,weight2_15;
Weight_MUX weight_mux2_0(.Weight_0(Wgt_2_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_2_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight2_0));
Weight_MUX weight_mux2_1(.Weight_0(Wgt_2_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_1));
Weight_MUX weight_mux2_2(.Weight_0(Wgt_2_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_2));
Weight_MUX weight_mux2_3(.Weight_0(Wgt_2_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_3));
Weight_MUX weight_mux2_4(.Weight_0(Wgt_2_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_4));
Weight_MUX weight_mux2_5(.Weight_0(Wgt_2_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_5));
Weight_MUX weight_mux2_6(.Weight_0(Wgt_2_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_6));
Weight_MUX weight_mux2_7(.Weight_0(Wgt_2_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_7));
Weight_MUX weight_mux2_8(.Weight_0(Wgt_2_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_8));
Weight_MUX weight_mux2_9(.Weight_0(Wgt_2_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_9));
Weight_MUX weight_mux2_10(.Weight_0(Wgt_2_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_10));
Weight_MUX weight_mux2_11(.Weight_0(Wgt_2_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_11));
Weight_MUX weight_mux2_12(.Weight_0(Wgt_2_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_12));
Weight_MUX weight_mux2_13(.Weight_0(Wgt_2_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_13));
Weight_MUX weight_mux2_14(.Weight_0(Wgt_2_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_14));
Weight_MUX weight_mux2_15(.Weight_0(Wgt_2_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_2_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_2_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_2_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_2_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_2_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_2_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_2_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_2_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_2_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_2_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_2_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_2_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_2_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_2_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_2_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_2_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_2_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_2_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_2_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_2_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_2_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_2_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_2_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_2_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_2_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_2_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_2_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_2_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_2_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_2_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_2_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_2_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_2_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_2_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_2_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_2_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_2_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_2_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_2_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_2_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_2_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_2_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_2_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_2_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_2_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_2_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_2_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_2_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight2_15));
wire [25:0] out_n2;
Neuron neuron_2(.Weight_0(weight2_0),.Weight_1(weight2_1),.Weight_2(weight2_2),.Weight_3(weight2_3),.Weight_4(weight2_4),.Weight_5(weight2_5),.Weight_6(weight2_6),.Weight_7(weight2_7),.Weight_8(weight2_8),.Weight_9(weight2_9),.Weight_10(weight2_10),.Weight_11(weight2_11),.Weight_12(weight2_12),.Weight_13(weight2_13),.Weight_14(weight2_14),.Weight_15(weight2_15),.Pixel_0(pixel2_0),.Pixel_1(pixel2_1),.Pixel_2(pixel2_2),.Pixel_3(pixel2_3),.Pixel_4(pixel2_4),.Pixel_5(pixel2_5),.Pixel_6(pixel2_6),.Pixel_7(pixel2_7),.Pixel_8(pixel2_8),.Pixel_9(pixel2_9),.Pixel_10(pixel2_10),.Pixel_11(pixel2_11),.Pixel_12(pixel2_12),.Pixel_13(pixel2_13),.Pixel_14(pixel2_14),.Pixel_15(pixel2_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n2));

// neuron_3
wire [`PIX_WIDTH-1:0] pixel3_0,pixel3_1,pixel3_2,pixel3_3,pixel3_4,pixel3_5,pixel3_6,pixel3_7,pixel3_8,pixel3_9,pixel3_10,pixel3_11,pixel3_12,pixel3_13,pixel3_14,pixel3_15;
Pixel_MUX pixel_mux3_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel3_0));
Pixel_MUX pixel_mux3_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_1));
Pixel_MUX pixel_mux3_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_2));
Pixel_MUX pixel_mux3_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_3));
Pixel_MUX pixel_mux3_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_4));
Pixel_MUX pixel_mux3_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_5));
Pixel_MUX pixel_mux3_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_6));
Pixel_MUX pixel_mux3_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_7));
Pixel_MUX pixel_mux3_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_8));
Pixel_MUX pixel_mux3_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_9));
Pixel_MUX pixel_mux3_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_10));
Pixel_MUX pixel_mux3_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_11));
Pixel_MUX pixel_mux3_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_12));
Pixel_MUX pixel_mux3_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_13));
Pixel_MUX pixel_mux3_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_14));
Pixel_MUX pixel_mux3_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel3_15));
wire [`WGT_WIDTH-1:0] weight3_0,weight3_1,weight3_2,weight3_3,weight3_4,weight3_5,weight3_6,weight3_7,weight3_8,weight3_9,weight3_10,weight3_11,weight3_12,weight3_13,weight3_14,weight3_15;
Weight_MUX weight_mux3_0(.Weight_0(Wgt_3_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_3_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight3_0));
Weight_MUX weight_mux3_1(.Weight_0(Wgt_3_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_1));
Weight_MUX weight_mux3_2(.Weight_0(Wgt_3_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_2));
Weight_MUX weight_mux3_3(.Weight_0(Wgt_3_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_3));
Weight_MUX weight_mux3_4(.Weight_0(Wgt_3_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_4));
Weight_MUX weight_mux3_5(.Weight_0(Wgt_3_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_5));
Weight_MUX weight_mux3_6(.Weight_0(Wgt_3_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_6));
Weight_MUX weight_mux3_7(.Weight_0(Wgt_3_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_7));
Weight_MUX weight_mux3_8(.Weight_0(Wgt_3_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_8));
Weight_MUX weight_mux3_9(.Weight_0(Wgt_3_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_9));
Weight_MUX weight_mux3_10(.Weight_0(Wgt_3_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_10));
Weight_MUX weight_mux3_11(.Weight_0(Wgt_3_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_11));
Weight_MUX weight_mux3_12(.Weight_0(Wgt_3_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_12));
Weight_MUX weight_mux3_13(.Weight_0(Wgt_3_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_13));
Weight_MUX weight_mux3_14(.Weight_0(Wgt_3_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_14));
Weight_MUX weight_mux3_15(.Weight_0(Wgt_3_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_3_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_3_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_3_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_3_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_3_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_3_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_3_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_3_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_3_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_3_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_3_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_3_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_3_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_3_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_3_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_3_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_3_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_3_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_3_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_3_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_3_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_3_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_3_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_3_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_3_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_3_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_3_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_3_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_3_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_3_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_3_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_3_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_3_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_3_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_3_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_3_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_3_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_3_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_3_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_3_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_3_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_3_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_3_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_3_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_3_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_3_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_3_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_3_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight3_15));
wire [25:0] out_n3;
Neuron neuron_3(.Weight_0(weight3_0),.Weight_1(weight3_1),.Weight_2(weight3_2),.Weight_3(weight3_3),.Weight_4(weight3_4),.Weight_5(weight3_5),.Weight_6(weight3_6),.Weight_7(weight3_7),.Weight_8(weight3_8),.Weight_9(weight3_9),.Weight_10(weight3_10),.Weight_11(weight3_11),.Weight_12(weight3_12),.Weight_13(weight3_13),.Weight_14(weight3_14),.Weight_15(weight3_15),.Pixel_0(pixel3_0),.Pixel_1(pixel3_1),.Pixel_2(pixel3_2),.Pixel_3(pixel3_3),.Pixel_4(pixel3_4),.Pixel_5(pixel3_5),.Pixel_6(pixel3_6),.Pixel_7(pixel3_7),.Pixel_8(pixel3_8),.Pixel_9(pixel3_9),.Pixel_10(pixel3_10),.Pixel_11(pixel3_11),.Pixel_12(pixel3_12),.Pixel_13(pixel3_13),.Pixel_14(pixel3_14),.Pixel_15(pixel3_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n3));

// neuron_4
wire [`PIX_WIDTH-1:0] pixel4_0,pixel4_1,pixel4_2,pixel4_3,pixel4_4,pixel4_5,pixel4_6,pixel4_7,pixel4_8,pixel4_9,pixel4_10,pixel4_11,pixel4_12,pixel4_13,pixel4_14,pixel4_15;
Pixel_MUX pixel_mux4_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel4_0));
Pixel_MUX pixel_mux4_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_1));
Pixel_MUX pixel_mux4_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_2));
Pixel_MUX pixel_mux4_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_3));
Pixel_MUX pixel_mux4_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_4));
Pixel_MUX pixel_mux4_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_5));
Pixel_MUX pixel_mux4_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_6));
Pixel_MUX pixel_mux4_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_7));
Pixel_MUX pixel_mux4_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_8));
Pixel_MUX pixel_mux4_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_9));
Pixel_MUX pixel_mux4_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_10));
Pixel_MUX pixel_mux4_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_11));
Pixel_MUX pixel_mux4_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_12));
Pixel_MUX pixel_mux4_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_13));
Pixel_MUX pixel_mux4_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_14));
Pixel_MUX pixel_mux4_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel4_15));
wire [`WGT_WIDTH-1:0] weight4_0,weight4_1,weight4_2,weight4_3,weight4_4,weight4_5,weight4_6,weight4_7,weight4_8,weight4_9,weight4_10,weight4_11,weight4_12,weight4_13,weight4_14,weight4_15;
Weight_MUX weight_mux4_0(.Weight_0(Wgt_4_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_4_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight4_0));
Weight_MUX weight_mux4_1(.Weight_0(Wgt_4_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_1));
Weight_MUX weight_mux4_2(.Weight_0(Wgt_4_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_2));
Weight_MUX weight_mux4_3(.Weight_0(Wgt_4_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_3));
Weight_MUX weight_mux4_4(.Weight_0(Wgt_4_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_4));
Weight_MUX weight_mux4_5(.Weight_0(Wgt_4_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_5));
Weight_MUX weight_mux4_6(.Weight_0(Wgt_4_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_6));
Weight_MUX weight_mux4_7(.Weight_0(Wgt_4_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_7));
Weight_MUX weight_mux4_8(.Weight_0(Wgt_4_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_8));
Weight_MUX weight_mux4_9(.Weight_0(Wgt_4_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_9));
Weight_MUX weight_mux4_10(.Weight_0(Wgt_4_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_10));
Weight_MUX weight_mux4_11(.Weight_0(Wgt_4_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_11));
Weight_MUX weight_mux4_12(.Weight_0(Wgt_4_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_12));
Weight_MUX weight_mux4_13(.Weight_0(Wgt_4_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_13));
Weight_MUX weight_mux4_14(.Weight_0(Wgt_4_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_14));
Weight_MUX weight_mux4_15(.Weight_0(Wgt_4_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_4_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_4_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_4_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_4_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_4_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_4_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_4_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_4_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_4_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_4_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_4_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_4_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_4_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_4_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_4_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_4_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_4_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_4_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_4_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_4_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_4_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_4_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_4_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_4_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_4_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_4_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_4_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_4_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_4_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_4_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_4_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_4_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_4_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_4_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_4_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_4_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_4_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_4_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_4_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_4_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_4_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_4_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_4_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_4_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_4_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_4_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_4_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_4_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight4_15));
wire [25:0] out_n4;
Neuron neuron_4(.Weight_0(weight4_0),.Weight_1(weight4_1),.Weight_2(weight4_2),.Weight_3(weight4_3),.Weight_4(weight4_4),.Weight_5(weight4_5),.Weight_6(weight4_6),.Weight_7(weight4_7),.Weight_8(weight4_8),.Weight_9(weight4_9),.Weight_10(weight4_10),.Weight_11(weight4_11),.Weight_12(weight4_12),.Weight_13(weight4_13),.Weight_14(weight4_14),.Weight_15(weight4_15),.Pixel_0(pixel4_0),.Pixel_1(pixel4_1),.Pixel_2(pixel4_2),.Pixel_3(pixel4_3),.Pixel_4(pixel4_4),.Pixel_5(pixel4_5),.Pixel_6(pixel4_6),.Pixel_7(pixel4_7),.Pixel_8(pixel4_8),.Pixel_9(pixel4_9),.Pixel_10(pixel4_10),.Pixel_11(pixel4_11),.Pixel_12(pixel4_12),.Pixel_13(pixel4_13),.Pixel_14(pixel4_14),.Pixel_15(pixel4_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n4));

// neuron_5
wire [`PIX_WIDTH-1:0] pixel5_0,pixel5_1,pixel5_2,pixel5_3,pixel5_4,pixel5_5,pixel5_6,pixel5_7,pixel5_8,pixel5_9,pixel5_10,pixel5_11,pixel5_12,pixel5_13,pixel5_14,pixel5_15;
Pixel_MUX pixel_mux5_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel5_0));
Pixel_MUX pixel_mux5_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_1));
Pixel_MUX pixel_mux5_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_2));
Pixel_MUX pixel_mux5_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_3));
Pixel_MUX pixel_mux5_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_4));
Pixel_MUX pixel_mux5_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_5));
Pixel_MUX pixel_mux5_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_6));
Pixel_MUX pixel_mux5_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_7));
Pixel_MUX pixel_mux5_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_8));
Pixel_MUX pixel_mux5_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_9));
Pixel_MUX pixel_mux5_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_10));
Pixel_MUX pixel_mux5_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_11));
Pixel_MUX pixel_mux5_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_12));
Pixel_MUX pixel_mux5_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_13));
Pixel_MUX pixel_mux5_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_14));
Pixel_MUX pixel_mux5_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel5_15));
wire [`WGT_WIDTH-1:0] weight5_0,weight5_1,weight5_2,weight5_3,weight5_4,weight5_5,weight5_6,weight5_7,weight5_8,weight5_9,weight5_10,weight5_11,weight5_12,weight5_13,weight5_14,weight5_15;
Weight_MUX weight_mux5_0(.Weight_0(Wgt_5_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_5_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight5_0));
Weight_MUX weight_mux5_1(.Weight_0(Wgt_5_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_1));
Weight_MUX weight_mux5_2(.Weight_0(Wgt_5_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_2));
Weight_MUX weight_mux5_3(.Weight_0(Wgt_5_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_3));
Weight_MUX weight_mux5_4(.Weight_0(Wgt_5_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_4));
Weight_MUX weight_mux5_5(.Weight_0(Wgt_5_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_5));
Weight_MUX weight_mux5_6(.Weight_0(Wgt_5_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_6));
Weight_MUX weight_mux5_7(.Weight_0(Wgt_5_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_7));
Weight_MUX weight_mux5_8(.Weight_0(Wgt_5_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_8));
Weight_MUX weight_mux5_9(.Weight_0(Wgt_5_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_9));
Weight_MUX weight_mux5_10(.Weight_0(Wgt_5_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_10));
Weight_MUX weight_mux5_11(.Weight_0(Wgt_5_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_11));
Weight_MUX weight_mux5_12(.Weight_0(Wgt_5_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_12));
Weight_MUX weight_mux5_13(.Weight_0(Wgt_5_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_13));
Weight_MUX weight_mux5_14(.Weight_0(Wgt_5_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_14));
Weight_MUX weight_mux5_15(.Weight_0(Wgt_5_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_5_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_5_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_5_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_5_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_5_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_5_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_5_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_5_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_5_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_5_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_5_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_5_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_5_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_5_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_5_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_5_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_5_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_5_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_5_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_5_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_5_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_5_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_5_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_5_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_5_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_5_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_5_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_5_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_5_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_5_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_5_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_5_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_5_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_5_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_5_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_5_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_5_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_5_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_5_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_5_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_5_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_5_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_5_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_5_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_5_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_5_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_5_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_5_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight5_15));
wire [25:0] out_n5;
Neuron neuron_5(.Weight_0(weight5_0),.Weight_1(weight5_1),.Weight_2(weight5_2),.Weight_3(weight5_3),.Weight_4(weight5_4),.Weight_5(weight5_5),.Weight_6(weight5_6),.Weight_7(weight5_7),.Weight_8(weight5_8),.Weight_9(weight5_9),.Weight_10(weight5_10),.Weight_11(weight5_11),.Weight_12(weight5_12),.Weight_13(weight5_13),.Weight_14(weight5_14),.Weight_15(weight5_15),.Pixel_0(pixel5_0),.Pixel_1(pixel5_1),.Pixel_2(pixel5_2),.Pixel_3(pixel5_3),.Pixel_4(pixel5_4),.Pixel_5(pixel5_5),.Pixel_6(pixel5_6),.Pixel_7(pixel5_7),.Pixel_8(pixel5_8),.Pixel_9(pixel5_9),.Pixel_10(pixel5_10),.Pixel_11(pixel5_11),.Pixel_12(pixel5_12),.Pixel_13(pixel5_13),.Pixel_14(pixel5_14),.Pixel_15(pixel5_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n5));

// neuron_6
wire [`PIX_WIDTH-1:0] pixel6_0,pixel6_1,pixel6_2,pixel6_3,pixel6_4,pixel6_5,pixel6_6,pixel6_7,pixel6_8,pixel6_9,pixel6_10,pixel6_11,pixel6_12,pixel6_13,pixel6_14,pixel6_15;
Pixel_MUX pixel_mux6_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel6_0));
Pixel_MUX pixel_mux6_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_1));
Pixel_MUX pixel_mux6_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_2));
Pixel_MUX pixel_mux6_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_3));
Pixel_MUX pixel_mux6_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_4));
Pixel_MUX pixel_mux6_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_5));
Pixel_MUX pixel_mux6_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_6));
Pixel_MUX pixel_mux6_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_7));
Pixel_MUX pixel_mux6_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_8));
Pixel_MUX pixel_mux6_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_9));
Pixel_MUX pixel_mux6_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_10));
Pixel_MUX pixel_mux6_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_11));
Pixel_MUX pixel_mux6_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_12));
Pixel_MUX pixel_mux6_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_13));
Pixel_MUX pixel_mux6_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_14));
Pixel_MUX pixel_mux6_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel6_15));
wire [`WGT_WIDTH-1:0] weight6_0,weight6_1,weight6_2,weight6_3,weight6_4,weight6_5,weight6_6,weight6_7,weight6_8,weight6_9,weight6_10,weight6_11,weight6_12,weight6_13,weight6_14,weight6_15;
Weight_MUX weight_mux6_0(.Weight_0(Wgt_6_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_6_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight6_0));
Weight_MUX weight_mux6_1(.Weight_0(Wgt_6_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_1));
Weight_MUX weight_mux6_2(.Weight_0(Wgt_6_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_2));
Weight_MUX weight_mux6_3(.Weight_0(Wgt_6_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_3));
Weight_MUX weight_mux6_4(.Weight_0(Wgt_6_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_4));
Weight_MUX weight_mux6_5(.Weight_0(Wgt_6_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_5));
Weight_MUX weight_mux6_6(.Weight_0(Wgt_6_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_6));
Weight_MUX weight_mux6_7(.Weight_0(Wgt_6_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_7));
Weight_MUX weight_mux6_8(.Weight_0(Wgt_6_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_8));
Weight_MUX weight_mux6_9(.Weight_0(Wgt_6_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_9));
Weight_MUX weight_mux6_10(.Weight_0(Wgt_6_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_10));
Weight_MUX weight_mux6_11(.Weight_0(Wgt_6_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_11));
Weight_MUX weight_mux6_12(.Weight_0(Wgt_6_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_12));
Weight_MUX weight_mux6_13(.Weight_0(Wgt_6_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_13));
Weight_MUX weight_mux6_14(.Weight_0(Wgt_6_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_14));
Weight_MUX weight_mux6_15(.Weight_0(Wgt_6_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_6_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_6_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_6_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_6_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_6_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_6_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_6_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_6_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_6_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_6_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_6_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_6_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_6_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_6_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_6_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_6_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_6_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_6_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_6_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_6_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_6_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_6_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_6_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_6_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_6_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_6_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_6_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_6_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_6_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_6_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_6_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_6_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_6_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_6_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_6_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_6_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_6_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_6_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_6_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_6_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_6_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_6_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_6_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_6_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_6_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_6_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_6_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_6_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight6_15));
wire [25:0] out_n6;
Neuron neuron_6(.Weight_0(weight6_0),.Weight_1(weight6_1),.Weight_2(weight6_2),.Weight_3(weight6_3),.Weight_4(weight6_4),.Weight_5(weight6_5),.Weight_6(weight6_6),.Weight_7(weight6_7),.Weight_8(weight6_8),.Weight_9(weight6_9),.Weight_10(weight6_10),.Weight_11(weight6_11),.Weight_12(weight6_12),.Weight_13(weight6_13),.Weight_14(weight6_14),.Weight_15(weight6_15),.Pixel_0(pixel6_0),.Pixel_1(pixel6_1),.Pixel_2(pixel6_2),.Pixel_3(pixel6_3),.Pixel_4(pixel6_4),.Pixel_5(pixel6_5),.Pixel_6(pixel6_6),.Pixel_7(pixel6_7),.Pixel_8(pixel6_8),.Pixel_9(pixel6_9),.Pixel_10(pixel6_10),.Pixel_11(pixel6_11),.Pixel_12(pixel6_12),.Pixel_13(pixel6_13),.Pixel_14(pixel6_14),.Pixel_15(pixel6_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n6));

// neuron_7
wire [`PIX_WIDTH-1:0] pixel7_0,pixel7_1,pixel7_2,pixel7_3,pixel7_4,pixel7_5,pixel7_6,pixel7_7,pixel7_8,pixel7_9,pixel7_10,pixel7_11,pixel7_12,pixel7_13,pixel7_14,pixel7_15;
Pixel_MUX pixel_mux7_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel7_0));
Pixel_MUX pixel_mux7_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_1));
Pixel_MUX pixel_mux7_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_2));
Pixel_MUX pixel_mux7_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_3));
Pixel_MUX pixel_mux7_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_4));
Pixel_MUX pixel_mux7_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_5));
Pixel_MUX pixel_mux7_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_6));
Pixel_MUX pixel_mux7_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_7));
Pixel_MUX pixel_mux7_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_8));
Pixel_MUX pixel_mux7_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_9));
Pixel_MUX pixel_mux7_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_10));
Pixel_MUX pixel_mux7_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_11));
Pixel_MUX pixel_mux7_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_12));
Pixel_MUX pixel_mux7_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_13));
Pixel_MUX pixel_mux7_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_14));
Pixel_MUX pixel_mux7_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel7_15));
wire [`WGT_WIDTH-1:0] weight7_0,weight7_1,weight7_2,weight7_3,weight7_4,weight7_5,weight7_6,weight7_7,weight7_8,weight7_9,weight7_10,weight7_11,weight7_12,weight7_13,weight7_14,weight7_15;
Weight_MUX weight_mux7_0(.Weight_0(Wgt_7_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_7_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight7_0));
Weight_MUX weight_mux7_1(.Weight_0(Wgt_7_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_1));
Weight_MUX weight_mux7_2(.Weight_0(Wgt_7_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_2));
Weight_MUX weight_mux7_3(.Weight_0(Wgt_7_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_3));
Weight_MUX weight_mux7_4(.Weight_0(Wgt_7_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_4));
Weight_MUX weight_mux7_5(.Weight_0(Wgt_7_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_5));
Weight_MUX weight_mux7_6(.Weight_0(Wgt_7_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_6));
Weight_MUX weight_mux7_7(.Weight_0(Wgt_7_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_7));
Weight_MUX weight_mux7_8(.Weight_0(Wgt_7_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_8));
Weight_MUX weight_mux7_9(.Weight_0(Wgt_7_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_9));
Weight_MUX weight_mux7_10(.Weight_0(Wgt_7_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_10));
Weight_MUX weight_mux7_11(.Weight_0(Wgt_7_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_11));
Weight_MUX weight_mux7_12(.Weight_0(Wgt_7_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_12));
Weight_MUX weight_mux7_13(.Weight_0(Wgt_7_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_13));
Weight_MUX weight_mux7_14(.Weight_0(Wgt_7_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_14));
Weight_MUX weight_mux7_15(.Weight_0(Wgt_7_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_7_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_7_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_7_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_7_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_7_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_7_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_7_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_7_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_7_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_7_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_7_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_7_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_7_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_7_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_7_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_7_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_7_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_7_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_7_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_7_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_7_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_7_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_7_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_7_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_7_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_7_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_7_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_7_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_7_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_7_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_7_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_7_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_7_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_7_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_7_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_7_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_7_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_7_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_7_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_7_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_7_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_7_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_7_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_7_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_7_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_7_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_7_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_7_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight7_15));
wire [25:0] out_n7;
Neuron neuron_7(.Weight_0(weight7_0),.Weight_1(weight7_1),.Weight_2(weight7_2),.Weight_3(weight7_3),.Weight_4(weight7_4),.Weight_5(weight7_5),.Weight_6(weight7_6),.Weight_7(weight7_7),.Weight_8(weight7_8),.Weight_9(weight7_9),.Weight_10(weight7_10),.Weight_11(weight7_11),.Weight_12(weight7_12),.Weight_13(weight7_13),.Weight_14(weight7_14),.Weight_15(weight7_15),.Pixel_0(pixel7_0),.Pixel_1(pixel7_1),.Pixel_2(pixel7_2),.Pixel_3(pixel7_3),.Pixel_4(pixel7_4),.Pixel_5(pixel7_5),.Pixel_6(pixel7_6),.Pixel_7(pixel7_7),.Pixel_8(pixel7_8),.Pixel_9(pixel7_9),.Pixel_10(pixel7_10),.Pixel_11(pixel7_11),.Pixel_12(pixel7_12),.Pixel_13(pixel7_13),.Pixel_14(pixel7_14),.Pixel_15(pixel7_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n7));

// neuron_8
wire [`PIX_WIDTH-1:0] pixel8_0,pixel8_1,pixel8_2,pixel8_3,pixel8_4,pixel8_5,pixel8_6,pixel8_7,pixel8_8,pixel8_9,pixel8_10,pixel8_11,pixel8_12,pixel8_13,pixel8_14,pixel8_15;
Pixel_MUX pixel_mux8_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel8_0));
Pixel_MUX pixel_mux8_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_1));
Pixel_MUX pixel_mux8_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_2));
Pixel_MUX pixel_mux8_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_3));
Pixel_MUX pixel_mux8_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_4));
Pixel_MUX pixel_mux8_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_5));
Pixel_MUX pixel_mux8_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_6));
Pixel_MUX pixel_mux8_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_7));
Pixel_MUX pixel_mux8_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_8));
Pixel_MUX pixel_mux8_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_9));
Pixel_MUX pixel_mux8_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_10));
Pixel_MUX pixel_mux8_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_11));
Pixel_MUX pixel_mux8_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_12));
Pixel_MUX pixel_mux8_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_13));
Pixel_MUX pixel_mux8_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_14));
Pixel_MUX pixel_mux8_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel8_15));
wire [`WGT_WIDTH-1:0] weight8_0,weight8_1,weight8_2,weight8_3,weight8_4,weight8_5,weight8_6,weight8_7,weight8_8,weight8_9,weight8_10,weight8_11,weight8_12,weight8_13,weight8_14,weight8_15;
Weight_MUX weight_mux8_0(.Weight_0(Wgt_8_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_8_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight8_0));
Weight_MUX weight_mux8_1(.Weight_0(Wgt_8_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_1));
Weight_MUX weight_mux8_2(.Weight_0(Wgt_8_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_2));
Weight_MUX weight_mux8_3(.Weight_0(Wgt_8_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_3));
Weight_MUX weight_mux8_4(.Weight_0(Wgt_8_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_4));
Weight_MUX weight_mux8_5(.Weight_0(Wgt_8_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_5));
Weight_MUX weight_mux8_6(.Weight_0(Wgt_8_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_6));
Weight_MUX weight_mux8_7(.Weight_0(Wgt_8_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_7));
Weight_MUX weight_mux8_8(.Weight_0(Wgt_8_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_8));
Weight_MUX weight_mux8_9(.Weight_0(Wgt_8_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_9));
Weight_MUX weight_mux8_10(.Weight_0(Wgt_8_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_10));
Weight_MUX weight_mux8_11(.Weight_0(Wgt_8_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_11));
Weight_MUX weight_mux8_12(.Weight_0(Wgt_8_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_12));
Weight_MUX weight_mux8_13(.Weight_0(Wgt_8_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_13));
Weight_MUX weight_mux8_14(.Weight_0(Wgt_8_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_14));
Weight_MUX weight_mux8_15(.Weight_0(Wgt_8_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_8_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_8_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_8_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_8_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_8_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_8_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_8_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_8_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_8_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_8_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_8_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_8_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_8_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_8_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_8_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_8_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_8_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_8_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_8_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_8_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_8_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_8_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_8_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_8_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_8_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_8_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_8_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_8_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_8_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_8_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_8_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_8_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_8_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_8_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_8_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_8_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_8_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_8_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_8_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_8_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_8_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_8_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_8_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_8_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_8_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_8_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_8_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_8_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight8_15));
wire [25:0] out_n8;
Neuron neuron_8(.Weight_0(weight8_0),.Weight_1(weight8_1),.Weight_2(weight8_2),.Weight_3(weight8_3),.Weight_4(weight8_4),.Weight_5(weight8_5),.Weight_6(weight8_6),.Weight_7(weight8_7),.Weight_8(weight8_8),.Weight_9(weight8_9),.Weight_10(weight8_10),.Weight_11(weight8_11),.Weight_12(weight8_12),.Weight_13(weight8_13),.Weight_14(weight8_14),.Weight_15(weight8_15),.Pixel_0(pixel8_0),.Pixel_1(pixel8_1),.Pixel_2(pixel8_2),.Pixel_3(pixel8_3),.Pixel_4(pixel8_4),.Pixel_5(pixel8_5),.Pixel_6(pixel8_6),.Pixel_7(pixel8_7),.Pixel_8(pixel8_8),.Pixel_9(pixel8_9),.Pixel_10(pixel8_10),.Pixel_11(pixel8_11),.Pixel_12(pixel8_12),.Pixel_13(pixel8_13),.Pixel_14(pixel8_14),.Pixel_15(pixel8_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n8));

// neuron_9
wire [`PIX_WIDTH-1:0] pixel9_0,pixel9_1,pixel9_2,pixel9_3,pixel9_4,pixel9_5,pixel9_6,pixel9_7,pixel9_8,pixel9_9,pixel9_10,pixel9_11,pixel9_12,pixel9_13,pixel9_14,pixel9_15;
Pixel_MUX pixel_mux9_0(.Pixel_0(Pixels[0]),.Pixel_1(Pixels[16]),.Pixel_2(Pixels[32]),.Pixel_3(Pixels[48]),.Pixel_4(Pixels[64]),.Pixel_5(Pixels[80]),.Pixel_6(Pixels[96]),.Pixel_7(Pixels[112]),.Pixel_8(Pixels[128]),.Pixel_9(Pixels[144]),.Pixel_10(Pixels[160]),.Pixel_11(Pixels[176]),.Pixel_12(Pixels[192]),.Pixel_13(Pixels[208]),.Pixel_14(Pixels[224]),.Pixel_15(Pixels[240]),.Pixel_16(Pixels[256]),.Pixel_17(Pixels[272]),.Pixel_18(Pixels[288]),.Pixel_19(Pixels[304]),.Pixel_20(Pixels[320]),.Pixel_21(Pixels[336]),.Pixel_22(Pixels[352]),.Pixel_23(Pixels[368]),.Pixel_24(Pixels[384]),.Pixel_25(Pixels[400]),.Pixel_26(Pixels[416]),.Pixel_27(Pixels[432]),.Pixel_28(Pixels[448]),.Pixel_29(Pixels[464]),.Pixel_30(Pixels[480]),.Pixel_31(Pixels[496]),.Pixel_32(Pixels[512]),.Pixel_33(Pixels[528]),.Pixel_34(Pixels[544]),.Pixel_35(Pixels[560]),.Pixel_36(Pixels[576]),.Pixel_37(Pixels[592]),.Pixel_38(Pixels[608]),.Pixel_39(Pixels[624]),.Pixel_40(Pixels[640]),.Pixel_41(Pixels[656]),.Pixel_42(Pixels[672]),.Pixel_43(Pixels[688]),.Pixel_44(Pixels[704]),.Pixel_45(Pixels[720]),.Pixel_46(Pixels[736]),.Pixel_47(Pixels[752]),.Pixel_48(Pixels[768]),.Pixel_49(Pixels[784]),.Pixel_Select(select_count),.Selected_Pixel(pixel9_0));
Pixel_MUX pixel_mux9_1(.Pixel_0(Pixels[1]),.Pixel_1(Pixels[17]),.Pixel_2(Pixels[33]),.Pixel_3(Pixels[49]),.Pixel_4(Pixels[65]),.Pixel_5(Pixels[81]),.Pixel_6(Pixels[97]),.Pixel_7(Pixels[113]),.Pixel_8(Pixels[129]),.Pixel_9(Pixels[145]),.Pixel_10(Pixels[161]),.Pixel_11(Pixels[177]),.Pixel_12(Pixels[193]),.Pixel_13(Pixels[209]),.Pixel_14(Pixels[225]),.Pixel_15(Pixels[241]),.Pixel_16(Pixels[257]),.Pixel_17(Pixels[273]),.Pixel_18(Pixels[289]),.Pixel_19(Pixels[305]),.Pixel_20(Pixels[321]),.Pixel_21(Pixels[337]),.Pixel_22(Pixels[353]),.Pixel_23(Pixels[369]),.Pixel_24(Pixels[385]),.Pixel_25(Pixels[401]),.Pixel_26(Pixels[417]),.Pixel_27(Pixels[433]),.Pixel_28(Pixels[449]),.Pixel_29(Pixels[465]),.Pixel_30(Pixels[481]),.Pixel_31(Pixels[497]),.Pixel_32(Pixels[513]),.Pixel_33(Pixels[529]),.Pixel_34(Pixels[545]),.Pixel_35(Pixels[561]),.Pixel_36(Pixels[577]),.Pixel_37(Pixels[593]),.Pixel_38(Pixels[609]),.Pixel_39(Pixels[625]),.Pixel_40(Pixels[641]),.Pixel_41(Pixels[657]),.Pixel_42(Pixels[673]),.Pixel_43(Pixels[689]),.Pixel_44(Pixels[705]),.Pixel_45(Pixels[721]),.Pixel_46(Pixels[737]),.Pixel_47(Pixels[753]),.Pixel_48(Pixels[769]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_1));
Pixel_MUX pixel_mux9_2(.Pixel_0(Pixels[2]),.Pixel_1(Pixels[18]),.Pixel_2(Pixels[34]),.Pixel_3(Pixels[50]),.Pixel_4(Pixels[66]),.Pixel_5(Pixels[82]),.Pixel_6(Pixels[98]),.Pixel_7(Pixels[114]),.Pixel_8(Pixels[130]),.Pixel_9(Pixels[146]),.Pixel_10(Pixels[162]),.Pixel_11(Pixels[178]),.Pixel_12(Pixels[194]),.Pixel_13(Pixels[210]),.Pixel_14(Pixels[226]),.Pixel_15(Pixels[242]),.Pixel_16(Pixels[258]),.Pixel_17(Pixels[274]),.Pixel_18(Pixels[290]),.Pixel_19(Pixels[306]),.Pixel_20(Pixels[322]),.Pixel_21(Pixels[338]),.Pixel_22(Pixels[354]),.Pixel_23(Pixels[370]),.Pixel_24(Pixels[386]),.Pixel_25(Pixels[402]),.Pixel_26(Pixels[418]),.Pixel_27(Pixels[434]),.Pixel_28(Pixels[450]),.Pixel_29(Pixels[466]),.Pixel_30(Pixels[482]),.Pixel_31(Pixels[498]),.Pixel_32(Pixels[514]),.Pixel_33(Pixels[530]),.Pixel_34(Pixels[546]),.Pixel_35(Pixels[562]),.Pixel_36(Pixels[578]),.Pixel_37(Pixels[594]),.Pixel_38(Pixels[610]),.Pixel_39(Pixels[626]),.Pixel_40(Pixels[642]),.Pixel_41(Pixels[658]),.Pixel_42(Pixels[674]),.Pixel_43(Pixels[690]),.Pixel_44(Pixels[706]),.Pixel_45(Pixels[722]),.Pixel_46(Pixels[738]),.Pixel_47(Pixels[754]),.Pixel_48(Pixels[770]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_2));
Pixel_MUX pixel_mux9_3(.Pixel_0(Pixels[3]),.Pixel_1(Pixels[19]),.Pixel_2(Pixels[35]),.Pixel_3(Pixels[51]),.Pixel_4(Pixels[67]),.Pixel_5(Pixels[83]),.Pixel_6(Pixels[99]),.Pixel_7(Pixels[115]),.Pixel_8(Pixels[131]),.Pixel_9(Pixels[147]),.Pixel_10(Pixels[163]),.Pixel_11(Pixels[179]),.Pixel_12(Pixels[195]),.Pixel_13(Pixels[211]),.Pixel_14(Pixels[227]),.Pixel_15(Pixels[243]),.Pixel_16(Pixels[259]),.Pixel_17(Pixels[275]),.Pixel_18(Pixels[291]),.Pixel_19(Pixels[307]),.Pixel_20(Pixels[323]),.Pixel_21(Pixels[339]),.Pixel_22(Pixels[355]),.Pixel_23(Pixels[371]),.Pixel_24(Pixels[387]),.Pixel_25(Pixels[403]),.Pixel_26(Pixels[419]),.Pixel_27(Pixels[435]),.Pixel_28(Pixels[451]),.Pixel_29(Pixels[467]),.Pixel_30(Pixels[483]),.Pixel_31(Pixels[499]),.Pixel_32(Pixels[515]),.Pixel_33(Pixels[531]),.Pixel_34(Pixels[547]),.Pixel_35(Pixels[563]),.Pixel_36(Pixels[579]),.Pixel_37(Pixels[595]),.Pixel_38(Pixels[611]),.Pixel_39(Pixels[627]),.Pixel_40(Pixels[643]),.Pixel_41(Pixels[659]),.Pixel_42(Pixels[675]),.Pixel_43(Pixels[691]),.Pixel_44(Pixels[707]),.Pixel_45(Pixels[723]),.Pixel_46(Pixels[739]),.Pixel_47(Pixels[755]),.Pixel_48(Pixels[771]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_3));
Pixel_MUX pixel_mux9_4(.Pixel_0(Pixels[4]),.Pixel_1(Pixels[20]),.Pixel_2(Pixels[36]),.Pixel_3(Pixels[52]),.Pixel_4(Pixels[68]),.Pixel_5(Pixels[84]),.Pixel_6(Pixels[100]),.Pixel_7(Pixels[116]),.Pixel_8(Pixels[132]),.Pixel_9(Pixels[148]),.Pixel_10(Pixels[164]),.Pixel_11(Pixels[180]),.Pixel_12(Pixels[196]),.Pixel_13(Pixels[212]),.Pixel_14(Pixels[228]),.Pixel_15(Pixels[244]),.Pixel_16(Pixels[260]),.Pixel_17(Pixels[276]),.Pixel_18(Pixels[292]),.Pixel_19(Pixels[308]),.Pixel_20(Pixels[324]),.Pixel_21(Pixels[340]),.Pixel_22(Pixels[356]),.Pixel_23(Pixels[372]),.Pixel_24(Pixels[388]),.Pixel_25(Pixels[404]),.Pixel_26(Pixels[420]),.Pixel_27(Pixels[436]),.Pixel_28(Pixels[452]),.Pixel_29(Pixels[468]),.Pixel_30(Pixels[484]),.Pixel_31(Pixels[500]),.Pixel_32(Pixels[516]),.Pixel_33(Pixels[532]),.Pixel_34(Pixels[548]),.Pixel_35(Pixels[564]),.Pixel_36(Pixels[580]),.Pixel_37(Pixels[596]),.Pixel_38(Pixels[612]),.Pixel_39(Pixels[628]),.Pixel_40(Pixels[644]),.Pixel_41(Pixels[660]),.Pixel_42(Pixels[676]),.Pixel_43(Pixels[692]),.Pixel_44(Pixels[708]),.Pixel_45(Pixels[724]),.Pixel_46(Pixels[740]),.Pixel_47(Pixels[756]),.Pixel_48(Pixels[772]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_4));
Pixel_MUX pixel_mux9_5(.Pixel_0(Pixels[5]),.Pixel_1(Pixels[21]),.Pixel_2(Pixels[37]),.Pixel_3(Pixels[53]),.Pixel_4(Pixels[69]),.Pixel_5(Pixels[85]),.Pixel_6(Pixels[101]),.Pixel_7(Pixels[117]),.Pixel_8(Pixels[133]),.Pixel_9(Pixels[149]),.Pixel_10(Pixels[165]),.Pixel_11(Pixels[181]),.Pixel_12(Pixels[197]),.Pixel_13(Pixels[213]),.Pixel_14(Pixels[229]),.Pixel_15(Pixels[245]),.Pixel_16(Pixels[261]),.Pixel_17(Pixels[277]),.Pixel_18(Pixels[293]),.Pixel_19(Pixels[309]),.Pixel_20(Pixels[325]),.Pixel_21(Pixels[341]),.Pixel_22(Pixels[357]),.Pixel_23(Pixels[373]),.Pixel_24(Pixels[389]),.Pixel_25(Pixels[405]),.Pixel_26(Pixels[421]),.Pixel_27(Pixels[437]),.Pixel_28(Pixels[453]),.Pixel_29(Pixels[469]),.Pixel_30(Pixels[485]),.Pixel_31(Pixels[501]),.Pixel_32(Pixels[517]),.Pixel_33(Pixels[533]),.Pixel_34(Pixels[549]),.Pixel_35(Pixels[565]),.Pixel_36(Pixels[581]),.Pixel_37(Pixels[597]),.Pixel_38(Pixels[613]),.Pixel_39(Pixels[629]),.Pixel_40(Pixels[645]),.Pixel_41(Pixels[661]),.Pixel_42(Pixels[677]),.Pixel_43(Pixels[693]),.Pixel_44(Pixels[709]),.Pixel_45(Pixels[725]),.Pixel_46(Pixels[741]),.Pixel_47(Pixels[757]),.Pixel_48(Pixels[773]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_5));
Pixel_MUX pixel_mux9_6(.Pixel_0(Pixels[6]),.Pixel_1(Pixels[22]),.Pixel_2(Pixels[38]),.Pixel_3(Pixels[54]),.Pixel_4(Pixels[70]),.Pixel_5(Pixels[86]),.Pixel_6(Pixels[102]),.Pixel_7(Pixels[118]),.Pixel_8(Pixels[134]),.Pixel_9(Pixels[150]),.Pixel_10(Pixels[166]),.Pixel_11(Pixels[182]),.Pixel_12(Pixels[198]),.Pixel_13(Pixels[214]),.Pixel_14(Pixels[230]),.Pixel_15(Pixels[246]),.Pixel_16(Pixels[262]),.Pixel_17(Pixels[278]),.Pixel_18(Pixels[294]),.Pixel_19(Pixels[310]),.Pixel_20(Pixels[326]),.Pixel_21(Pixels[342]),.Pixel_22(Pixels[358]),.Pixel_23(Pixels[374]),.Pixel_24(Pixels[390]),.Pixel_25(Pixels[406]),.Pixel_26(Pixels[422]),.Pixel_27(Pixels[438]),.Pixel_28(Pixels[454]),.Pixel_29(Pixels[470]),.Pixel_30(Pixels[486]),.Pixel_31(Pixels[502]),.Pixel_32(Pixels[518]),.Pixel_33(Pixels[534]),.Pixel_34(Pixels[550]),.Pixel_35(Pixels[566]),.Pixel_36(Pixels[582]),.Pixel_37(Pixels[598]),.Pixel_38(Pixels[614]),.Pixel_39(Pixels[630]),.Pixel_40(Pixels[646]),.Pixel_41(Pixels[662]),.Pixel_42(Pixels[678]),.Pixel_43(Pixels[694]),.Pixel_44(Pixels[710]),.Pixel_45(Pixels[726]),.Pixel_46(Pixels[742]),.Pixel_47(Pixels[758]),.Pixel_48(Pixels[774]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_6));
Pixel_MUX pixel_mux9_7(.Pixel_0(Pixels[7]),.Pixel_1(Pixels[23]),.Pixel_2(Pixels[39]),.Pixel_3(Pixels[55]),.Pixel_4(Pixels[71]),.Pixel_5(Pixels[87]),.Pixel_6(Pixels[103]),.Pixel_7(Pixels[119]),.Pixel_8(Pixels[135]),.Pixel_9(Pixels[151]),.Pixel_10(Pixels[167]),.Pixel_11(Pixels[183]),.Pixel_12(Pixels[199]),.Pixel_13(Pixels[215]),.Pixel_14(Pixels[231]),.Pixel_15(Pixels[247]),.Pixel_16(Pixels[263]),.Pixel_17(Pixels[279]),.Pixel_18(Pixels[295]),.Pixel_19(Pixels[311]),.Pixel_20(Pixels[327]),.Pixel_21(Pixels[343]),.Pixel_22(Pixels[359]),.Pixel_23(Pixels[375]),.Pixel_24(Pixels[391]),.Pixel_25(Pixels[407]),.Pixel_26(Pixels[423]),.Pixel_27(Pixels[439]),.Pixel_28(Pixels[455]),.Pixel_29(Pixels[471]),.Pixel_30(Pixels[487]),.Pixel_31(Pixels[503]),.Pixel_32(Pixels[519]),.Pixel_33(Pixels[535]),.Pixel_34(Pixels[551]),.Pixel_35(Pixels[567]),.Pixel_36(Pixels[583]),.Pixel_37(Pixels[599]),.Pixel_38(Pixels[615]),.Pixel_39(Pixels[631]),.Pixel_40(Pixels[647]),.Pixel_41(Pixels[663]),.Pixel_42(Pixels[679]),.Pixel_43(Pixels[695]),.Pixel_44(Pixels[711]),.Pixel_45(Pixels[727]),.Pixel_46(Pixels[743]),.Pixel_47(Pixels[759]),.Pixel_48(Pixels[775]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_7));
Pixel_MUX pixel_mux9_8(.Pixel_0(Pixels[8]),.Pixel_1(Pixels[24]),.Pixel_2(Pixels[40]),.Pixel_3(Pixels[56]),.Pixel_4(Pixels[72]),.Pixel_5(Pixels[88]),.Pixel_6(Pixels[104]),.Pixel_7(Pixels[120]),.Pixel_8(Pixels[136]),.Pixel_9(Pixels[152]),.Pixel_10(Pixels[168]),.Pixel_11(Pixels[184]),.Pixel_12(Pixels[200]),.Pixel_13(Pixels[216]),.Pixel_14(Pixels[232]),.Pixel_15(Pixels[248]),.Pixel_16(Pixels[264]),.Pixel_17(Pixels[280]),.Pixel_18(Pixels[296]),.Pixel_19(Pixels[312]),.Pixel_20(Pixels[328]),.Pixel_21(Pixels[344]),.Pixel_22(Pixels[360]),.Pixel_23(Pixels[376]),.Pixel_24(Pixels[392]),.Pixel_25(Pixels[408]),.Pixel_26(Pixels[424]),.Pixel_27(Pixels[440]),.Pixel_28(Pixels[456]),.Pixel_29(Pixels[472]),.Pixel_30(Pixels[488]),.Pixel_31(Pixels[504]),.Pixel_32(Pixels[520]),.Pixel_33(Pixels[536]),.Pixel_34(Pixels[552]),.Pixel_35(Pixels[568]),.Pixel_36(Pixels[584]),.Pixel_37(Pixels[600]),.Pixel_38(Pixels[616]),.Pixel_39(Pixels[632]),.Pixel_40(Pixels[648]),.Pixel_41(Pixels[664]),.Pixel_42(Pixels[680]),.Pixel_43(Pixels[696]),.Pixel_44(Pixels[712]),.Pixel_45(Pixels[728]),.Pixel_46(Pixels[744]),.Pixel_47(Pixels[760]),.Pixel_48(Pixels[776]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_8));
Pixel_MUX pixel_mux9_9(.Pixel_0(Pixels[9]),.Pixel_1(Pixels[25]),.Pixel_2(Pixels[41]),.Pixel_3(Pixels[57]),.Pixel_4(Pixels[73]),.Pixel_5(Pixels[89]),.Pixel_6(Pixels[105]),.Pixel_7(Pixels[121]),.Pixel_8(Pixels[137]),.Pixel_9(Pixels[153]),.Pixel_10(Pixels[169]),.Pixel_11(Pixels[185]),.Pixel_12(Pixels[201]),.Pixel_13(Pixels[217]),.Pixel_14(Pixels[233]),.Pixel_15(Pixels[249]),.Pixel_16(Pixels[265]),.Pixel_17(Pixels[281]),.Pixel_18(Pixels[297]),.Pixel_19(Pixels[313]),.Pixel_20(Pixels[329]),.Pixel_21(Pixels[345]),.Pixel_22(Pixels[361]),.Pixel_23(Pixels[377]),.Pixel_24(Pixels[393]),.Pixel_25(Pixels[409]),.Pixel_26(Pixels[425]),.Pixel_27(Pixels[441]),.Pixel_28(Pixels[457]),.Pixel_29(Pixels[473]),.Pixel_30(Pixels[489]),.Pixel_31(Pixels[505]),.Pixel_32(Pixels[521]),.Pixel_33(Pixels[537]),.Pixel_34(Pixels[553]),.Pixel_35(Pixels[569]),.Pixel_36(Pixels[585]),.Pixel_37(Pixels[601]),.Pixel_38(Pixels[617]),.Pixel_39(Pixels[633]),.Pixel_40(Pixels[649]),.Pixel_41(Pixels[665]),.Pixel_42(Pixels[681]),.Pixel_43(Pixels[697]),.Pixel_44(Pixels[713]),.Pixel_45(Pixels[729]),.Pixel_46(Pixels[745]),.Pixel_47(Pixels[761]),.Pixel_48(Pixels[777]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_9));
Pixel_MUX pixel_mux9_10(.Pixel_0(Pixels[10]),.Pixel_1(Pixels[26]),.Pixel_2(Pixels[42]),.Pixel_3(Pixels[58]),.Pixel_4(Pixels[74]),.Pixel_5(Pixels[90]),.Pixel_6(Pixels[106]),.Pixel_7(Pixels[122]),.Pixel_8(Pixels[138]),.Pixel_9(Pixels[154]),.Pixel_10(Pixels[170]),.Pixel_11(Pixels[186]),.Pixel_12(Pixels[202]),.Pixel_13(Pixels[218]),.Pixel_14(Pixels[234]),.Pixel_15(Pixels[250]),.Pixel_16(Pixels[266]),.Pixel_17(Pixels[282]),.Pixel_18(Pixels[298]),.Pixel_19(Pixels[314]),.Pixel_20(Pixels[330]),.Pixel_21(Pixels[346]),.Pixel_22(Pixels[362]),.Pixel_23(Pixels[378]),.Pixel_24(Pixels[394]),.Pixel_25(Pixels[410]),.Pixel_26(Pixels[426]),.Pixel_27(Pixels[442]),.Pixel_28(Pixels[458]),.Pixel_29(Pixels[474]),.Pixel_30(Pixels[490]),.Pixel_31(Pixels[506]),.Pixel_32(Pixels[522]),.Pixel_33(Pixels[538]),.Pixel_34(Pixels[554]),.Pixel_35(Pixels[570]),.Pixel_36(Pixels[586]),.Pixel_37(Pixels[602]),.Pixel_38(Pixels[618]),.Pixel_39(Pixels[634]),.Pixel_40(Pixels[650]),.Pixel_41(Pixels[666]),.Pixel_42(Pixels[682]),.Pixel_43(Pixels[698]),.Pixel_44(Pixels[714]),.Pixel_45(Pixels[730]),.Pixel_46(Pixels[746]),.Pixel_47(Pixels[762]),.Pixel_48(Pixels[778]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_10));
Pixel_MUX pixel_mux9_11(.Pixel_0(Pixels[11]),.Pixel_1(Pixels[27]),.Pixel_2(Pixels[43]),.Pixel_3(Pixels[59]),.Pixel_4(Pixels[75]),.Pixel_5(Pixels[91]),.Pixel_6(Pixels[107]),.Pixel_7(Pixels[123]),.Pixel_8(Pixels[139]),.Pixel_9(Pixels[155]),.Pixel_10(Pixels[171]),.Pixel_11(Pixels[187]),.Pixel_12(Pixels[203]),.Pixel_13(Pixels[219]),.Pixel_14(Pixels[235]),.Pixel_15(Pixels[251]),.Pixel_16(Pixels[267]),.Pixel_17(Pixels[283]),.Pixel_18(Pixels[299]),.Pixel_19(Pixels[315]),.Pixel_20(Pixels[331]),.Pixel_21(Pixels[347]),.Pixel_22(Pixels[363]),.Pixel_23(Pixels[379]),.Pixel_24(Pixels[395]),.Pixel_25(Pixels[411]),.Pixel_26(Pixels[427]),.Pixel_27(Pixels[443]),.Pixel_28(Pixels[459]),.Pixel_29(Pixels[475]),.Pixel_30(Pixels[491]),.Pixel_31(Pixels[507]),.Pixel_32(Pixels[523]),.Pixel_33(Pixels[539]),.Pixel_34(Pixels[555]),.Pixel_35(Pixels[571]),.Pixel_36(Pixels[587]),.Pixel_37(Pixels[603]),.Pixel_38(Pixels[619]),.Pixel_39(Pixels[635]),.Pixel_40(Pixels[651]),.Pixel_41(Pixels[667]),.Pixel_42(Pixels[683]),.Pixel_43(Pixels[699]),.Pixel_44(Pixels[715]),.Pixel_45(Pixels[731]),.Pixel_46(Pixels[747]),.Pixel_47(Pixels[763]),.Pixel_48(Pixels[779]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_11));
Pixel_MUX pixel_mux9_12(.Pixel_0(Pixels[12]),.Pixel_1(Pixels[28]),.Pixel_2(Pixels[44]),.Pixel_3(Pixels[60]),.Pixel_4(Pixels[76]),.Pixel_5(Pixels[92]),.Pixel_6(Pixels[108]),.Pixel_7(Pixels[124]),.Pixel_8(Pixels[140]),.Pixel_9(Pixels[156]),.Pixel_10(Pixels[172]),.Pixel_11(Pixels[188]),.Pixel_12(Pixels[204]),.Pixel_13(Pixels[220]),.Pixel_14(Pixels[236]),.Pixel_15(Pixels[252]),.Pixel_16(Pixels[268]),.Pixel_17(Pixels[284]),.Pixel_18(Pixels[300]),.Pixel_19(Pixels[316]),.Pixel_20(Pixels[332]),.Pixel_21(Pixels[348]),.Pixel_22(Pixels[364]),.Pixel_23(Pixels[380]),.Pixel_24(Pixels[396]),.Pixel_25(Pixels[412]),.Pixel_26(Pixels[428]),.Pixel_27(Pixels[444]),.Pixel_28(Pixels[460]),.Pixel_29(Pixels[476]),.Pixel_30(Pixels[492]),.Pixel_31(Pixels[508]),.Pixel_32(Pixels[524]),.Pixel_33(Pixels[540]),.Pixel_34(Pixels[556]),.Pixel_35(Pixels[572]),.Pixel_36(Pixels[588]),.Pixel_37(Pixels[604]),.Pixel_38(Pixels[620]),.Pixel_39(Pixels[636]),.Pixel_40(Pixels[652]),.Pixel_41(Pixels[668]),.Pixel_42(Pixels[684]),.Pixel_43(Pixels[700]),.Pixel_44(Pixels[716]),.Pixel_45(Pixels[732]),.Pixel_46(Pixels[748]),.Pixel_47(Pixels[764]),.Pixel_48(Pixels[780]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_12));
Pixel_MUX pixel_mux9_13(.Pixel_0(Pixels[13]),.Pixel_1(Pixels[29]),.Pixel_2(Pixels[45]),.Pixel_3(Pixels[61]),.Pixel_4(Pixels[77]),.Pixel_5(Pixels[93]),.Pixel_6(Pixels[109]),.Pixel_7(Pixels[125]),.Pixel_8(Pixels[141]),.Pixel_9(Pixels[157]),.Pixel_10(Pixels[173]),.Pixel_11(Pixels[189]),.Pixel_12(Pixels[205]),.Pixel_13(Pixels[221]),.Pixel_14(Pixels[237]),.Pixel_15(Pixels[253]),.Pixel_16(Pixels[269]),.Pixel_17(Pixels[285]),.Pixel_18(Pixels[301]),.Pixel_19(Pixels[317]),.Pixel_20(Pixels[333]),.Pixel_21(Pixels[349]),.Pixel_22(Pixels[365]),.Pixel_23(Pixels[381]),.Pixel_24(Pixels[397]),.Pixel_25(Pixels[413]),.Pixel_26(Pixels[429]),.Pixel_27(Pixels[445]),.Pixel_28(Pixels[461]),.Pixel_29(Pixels[477]),.Pixel_30(Pixels[493]),.Pixel_31(Pixels[509]),.Pixel_32(Pixels[525]),.Pixel_33(Pixels[541]),.Pixel_34(Pixels[557]),.Pixel_35(Pixels[573]),.Pixel_36(Pixels[589]),.Pixel_37(Pixels[605]),.Pixel_38(Pixels[621]),.Pixel_39(Pixels[637]),.Pixel_40(Pixels[653]),.Pixel_41(Pixels[669]),.Pixel_42(Pixels[685]),.Pixel_43(Pixels[701]),.Pixel_44(Pixels[717]),.Pixel_45(Pixels[733]),.Pixel_46(Pixels[749]),.Pixel_47(Pixels[765]),.Pixel_48(Pixels[781]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_13));
Pixel_MUX pixel_mux9_14(.Pixel_0(Pixels[14]),.Pixel_1(Pixels[30]),.Pixel_2(Pixels[46]),.Pixel_3(Pixels[62]),.Pixel_4(Pixels[78]),.Pixel_5(Pixels[94]),.Pixel_6(Pixels[110]),.Pixel_7(Pixels[126]),.Pixel_8(Pixels[142]),.Pixel_9(Pixels[158]),.Pixel_10(Pixels[174]),.Pixel_11(Pixels[190]),.Pixel_12(Pixels[206]),.Pixel_13(Pixels[222]),.Pixel_14(Pixels[238]),.Pixel_15(Pixels[254]),.Pixel_16(Pixels[270]),.Pixel_17(Pixels[286]),.Pixel_18(Pixels[302]),.Pixel_19(Pixels[318]),.Pixel_20(Pixels[334]),.Pixel_21(Pixels[350]),.Pixel_22(Pixels[366]),.Pixel_23(Pixels[382]),.Pixel_24(Pixels[398]),.Pixel_25(Pixels[414]),.Pixel_26(Pixels[430]),.Pixel_27(Pixels[446]),.Pixel_28(Pixels[462]),.Pixel_29(Pixels[478]),.Pixel_30(Pixels[494]),.Pixel_31(Pixels[510]),.Pixel_32(Pixels[526]),.Pixel_33(Pixels[542]),.Pixel_34(Pixels[558]),.Pixel_35(Pixels[574]),.Pixel_36(Pixels[590]),.Pixel_37(Pixels[606]),.Pixel_38(Pixels[622]),.Pixel_39(Pixels[638]),.Pixel_40(Pixels[654]),.Pixel_41(Pixels[670]),.Pixel_42(Pixels[686]),.Pixel_43(Pixels[702]),.Pixel_44(Pixels[718]),.Pixel_45(Pixels[734]),.Pixel_46(Pixels[750]),.Pixel_47(Pixels[766]),.Pixel_48(Pixels[782]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_14));
Pixel_MUX pixel_mux9_15(.Pixel_0(Pixels[15]),.Pixel_1(Pixels[31]),.Pixel_2(Pixels[47]),.Pixel_3(Pixels[63]),.Pixel_4(Pixels[79]),.Pixel_5(Pixels[95]),.Pixel_6(Pixels[111]),.Pixel_7(Pixels[127]),.Pixel_8(Pixels[143]),.Pixel_9(Pixels[159]),.Pixel_10(Pixels[175]),.Pixel_11(Pixels[191]),.Pixel_12(Pixels[207]),.Pixel_13(Pixels[223]),.Pixel_14(Pixels[239]),.Pixel_15(Pixels[255]),.Pixel_16(Pixels[271]),.Pixel_17(Pixels[287]),.Pixel_18(Pixels[303]),.Pixel_19(Pixels[319]),.Pixel_20(Pixels[335]),.Pixel_21(Pixels[351]),.Pixel_22(Pixels[367]),.Pixel_23(Pixels[383]),.Pixel_24(Pixels[399]),.Pixel_25(Pixels[415]),.Pixel_26(Pixels[431]),.Pixel_27(Pixels[447]),.Pixel_28(Pixels[463]),.Pixel_29(Pixels[479]),.Pixel_30(Pixels[495]),.Pixel_31(Pixels[511]),.Pixel_32(Pixels[527]),.Pixel_33(Pixels[543]),.Pixel_34(Pixels[559]),.Pixel_35(Pixels[575]),.Pixel_36(Pixels[591]),.Pixel_37(Pixels[607]),.Pixel_38(Pixels[623]),.Pixel_39(Pixels[639]),.Pixel_40(Pixels[655]),.Pixel_41(Pixels[671]),.Pixel_42(Pixels[687]),.Pixel_43(Pixels[703]),.Pixel_44(Pixels[719]),.Pixel_45(Pixels[735]),.Pixel_46(Pixels[751]),.Pixel_47(Pixels[767]),.Pixel_48(Pixels[783]),.Pixel_49(`PIX_WIDTH'b0),.Pixel_Select(select_count),.Selected_Pixel(pixel9_15));
wire [`WGT_WIDTH-1:0] weight9_0,weight9_1,weight9_2,weight9_3,weight9_4,weight9_5,weight9_6,weight9_7,weight9_8,weight9_9,weight9_10,weight9_11,weight9_12,weight9_13,weight9_14,weight9_15;
Weight_MUX weight_mux9_0(.Weight_0(Wgt_9_0[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_16[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_32[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_48[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_64[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_80[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_96[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_112[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_128[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_144[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_160[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_176[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_192[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_208[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_224[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_240[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_256[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_272[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_288[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_304[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_320[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_336[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_352[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_368[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_384[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_400[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_416[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_432[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_448[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_464[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_480[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_496[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_512[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_528[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_544[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_560[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_576[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_592[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_608[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_624[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_640[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_656[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_672[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_688[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_704[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_720[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_736[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_752[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_768[18:19-`WGT_WIDTH]),.Weight_49(Wgt_9_784[18:19-`WGT_WIDTH]),.Weight_Select(select_count),.Selected_Weight(weight9_0));
Weight_MUX weight_mux9_1(.Weight_0(Wgt_9_1[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_17[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_33[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_49[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_65[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_81[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_97[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_113[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_129[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_145[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_161[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_177[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_193[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_209[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_225[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_241[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_257[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_273[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_289[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_305[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_321[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_337[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_353[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_369[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_385[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_401[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_417[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_433[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_449[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_465[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_481[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_497[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_513[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_529[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_545[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_561[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_577[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_593[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_609[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_625[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_641[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_657[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_673[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_689[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_705[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_721[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_737[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_753[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_769[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_1));
Weight_MUX weight_mux9_2(.Weight_0(Wgt_9_2[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_18[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_34[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_50[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_66[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_82[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_98[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_114[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_130[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_146[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_162[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_178[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_194[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_210[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_226[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_242[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_258[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_274[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_290[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_306[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_322[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_338[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_354[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_370[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_386[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_402[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_418[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_434[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_450[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_466[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_482[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_498[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_514[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_530[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_546[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_562[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_578[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_594[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_610[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_626[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_642[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_658[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_674[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_690[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_706[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_722[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_738[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_754[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_770[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_2));
Weight_MUX weight_mux9_3(.Weight_0(Wgt_9_3[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_19[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_35[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_51[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_67[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_83[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_99[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_115[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_131[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_147[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_163[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_179[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_195[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_211[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_227[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_243[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_259[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_275[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_291[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_307[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_323[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_339[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_355[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_371[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_387[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_403[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_419[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_435[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_451[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_467[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_483[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_499[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_515[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_531[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_547[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_563[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_579[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_595[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_611[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_627[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_643[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_659[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_675[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_691[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_707[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_723[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_739[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_755[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_771[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_3));
Weight_MUX weight_mux9_4(.Weight_0(Wgt_9_4[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_20[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_36[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_52[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_68[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_84[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_100[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_116[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_132[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_148[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_164[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_180[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_196[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_212[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_228[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_244[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_260[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_276[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_292[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_308[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_324[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_340[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_356[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_372[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_388[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_404[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_420[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_436[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_452[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_468[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_484[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_500[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_516[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_532[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_548[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_564[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_580[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_596[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_612[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_628[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_644[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_660[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_676[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_692[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_708[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_724[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_740[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_756[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_772[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_4));
Weight_MUX weight_mux9_5(.Weight_0(Wgt_9_5[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_21[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_37[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_53[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_69[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_85[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_101[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_117[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_133[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_149[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_165[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_181[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_197[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_213[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_229[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_245[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_261[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_277[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_293[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_309[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_325[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_341[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_357[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_373[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_389[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_405[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_421[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_437[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_453[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_469[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_485[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_501[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_517[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_533[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_549[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_565[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_581[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_597[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_613[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_629[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_645[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_661[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_677[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_693[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_709[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_725[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_741[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_757[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_773[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_5));
Weight_MUX weight_mux9_6(.Weight_0(Wgt_9_6[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_22[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_38[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_54[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_70[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_86[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_102[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_118[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_134[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_150[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_166[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_182[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_198[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_214[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_230[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_246[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_262[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_278[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_294[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_310[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_326[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_342[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_358[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_374[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_390[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_406[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_422[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_438[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_454[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_470[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_486[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_502[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_518[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_534[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_550[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_566[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_582[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_598[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_614[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_630[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_646[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_662[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_678[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_694[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_710[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_726[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_742[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_758[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_774[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_6));
Weight_MUX weight_mux9_7(.Weight_0(Wgt_9_7[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_23[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_39[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_55[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_71[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_87[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_103[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_119[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_135[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_151[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_167[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_183[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_199[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_215[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_231[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_247[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_263[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_279[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_295[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_311[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_327[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_343[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_359[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_375[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_391[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_407[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_423[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_439[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_455[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_471[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_487[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_503[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_519[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_535[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_551[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_567[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_583[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_599[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_615[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_631[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_647[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_663[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_679[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_695[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_711[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_727[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_743[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_759[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_775[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_7));
Weight_MUX weight_mux9_8(.Weight_0(Wgt_9_8[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_24[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_40[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_56[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_72[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_88[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_104[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_120[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_136[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_152[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_168[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_184[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_200[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_216[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_232[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_248[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_264[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_280[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_296[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_312[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_328[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_344[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_360[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_376[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_392[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_408[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_424[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_440[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_456[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_472[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_488[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_504[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_520[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_536[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_552[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_568[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_584[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_600[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_616[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_632[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_648[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_664[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_680[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_696[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_712[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_728[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_744[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_760[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_776[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_8));
Weight_MUX weight_mux9_9(.Weight_0(Wgt_9_9[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_25[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_41[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_57[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_73[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_89[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_105[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_121[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_137[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_153[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_169[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_185[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_201[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_217[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_233[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_249[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_265[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_281[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_297[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_313[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_329[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_345[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_361[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_377[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_393[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_409[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_425[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_441[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_457[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_473[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_489[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_505[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_521[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_537[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_553[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_569[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_585[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_601[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_617[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_633[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_649[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_665[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_681[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_697[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_713[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_729[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_745[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_761[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_777[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_9));
Weight_MUX weight_mux9_10(.Weight_0(Wgt_9_10[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_26[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_42[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_58[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_74[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_90[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_106[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_122[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_138[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_154[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_170[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_186[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_202[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_218[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_234[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_250[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_266[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_282[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_298[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_314[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_330[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_346[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_362[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_378[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_394[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_410[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_426[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_442[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_458[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_474[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_490[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_506[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_522[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_538[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_554[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_570[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_586[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_602[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_618[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_634[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_650[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_666[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_682[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_698[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_714[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_730[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_746[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_762[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_778[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_10));
Weight_MUX weight_mux9_11(.Weight_0(Wgt_9_11[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_27[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_43[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_59[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_75[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_91[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_107[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_123[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_139[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_155[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_171[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_187[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_203[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_219[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_235[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_251[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_267[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_283[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_299[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_315[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_331[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_347[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_363[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_379[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_395[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_411[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_427[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_443[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_459[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_475[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_491[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_507[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_523[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_539[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_555[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_571[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_587[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_603[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_619[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_635[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_651[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_667[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_683[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_699[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_715[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_731[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_747[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_763[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_779[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_11));
Weight_MUX weight_mux9_12(.Weight_0(Wgt_9_12[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_28[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_44[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_60[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_76[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_92[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_108[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_124[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_140[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_156[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_172[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_188[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_204[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_220[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_236[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_252[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_268[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_284[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_300[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_316[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_332[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_348[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_364[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_380[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_396[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_412[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_428[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_444[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_460[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_476[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_492[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_508[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_524[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_540[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_556[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_572[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_588[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_604[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_620[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_636[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_652[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_668[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_684[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_700[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_716[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_732[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_748[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_764[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_780[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_12));
Weight_MUX weight_mux9_13(.Weight_0(Wgt_9_13[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_29[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_45[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_61[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_77[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_93[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_109[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_125[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_141[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_157[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_173[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_189[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_205[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_221[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_237[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_253[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_269[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_285[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_301[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_317[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_333[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_349[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_365[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_381[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_397[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_413[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_429[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_445[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_461[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_477[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_493[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_509[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_525[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_541[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_557[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_573[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_589[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_605[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_621[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_637[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_653[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_669[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_685[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_701[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_717[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_733[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_749[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_765[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_781[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_13));
Weight_MUX weight_mux9_14(.Weight_0(Wgt_9_14[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_30[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_46[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_62[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_78[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_94[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_110[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_126[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_142[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_158[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_174[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_190[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_206[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_222[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_238[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_254[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_270[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_286[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_302[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_318[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_334[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_350[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_366[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_382[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_398[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_414[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_430[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_446[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_462[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_478[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_494[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_510[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_526[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_542[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_558[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_574[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_590[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_606[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_622[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_638[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_654[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_670[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_686[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_702[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_718[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_734[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_750[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_766[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_782[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_14));
Weight_MUX weight_mux9_15(.Weight_0(Wgt_9_15[18:19-`WGT_WIDTH]),.Weight_1(Wgt_9_31[18:19-`WGT_WIDTH]),.Weight_2(Wgt_9_47[18:19-`WGT_WIDTH]),.Weight_3(Wgt_9_63[18:19-`WGT_WIDTH]),.Weight_4(Wgt_9_79[18:19-`WGT_WIDTH]),.Weight_5(Wgt_9_95[18:19-`WGT_WIDTH]),.Weight_6(Wgt_9_111[18:19-`WGT_WIDTH]),.Weight_7(Wgt_9_127[18:19-`WGT_WIDTH]),.Weight_8(Wgt_9_143[18:19-`WGT_WIDTH]),.Weight_9(Wgt_9_159[18:19-`WGT_WIDTH]),.Weight_10(Wgt_9_175[18:19-`WGT_WIDTH]),.Weight_11(Wgt_9_191[18:19-`WGT_WIDTH]),.Weight_12(Wgt_9_207[18:19-`WGT_WIDTH]),.Weight_13(Wgt_9_223[18:19-`WGT_WIDTH]),.Weight_14(Wgt_9_239[18:19-`WGT_WIDTH]),.Weight_15(Wgt_9_255[18:19-`WGT_WIDTH]),.Weight_16(Wgt_9_271[18:19-`WGT_WIDTH]),.Weight_17(Wgt_9_287[18:19-`WGT_WIDTH]),.Weight_18(Wgt_9_303[18:19-`WGT_WIDTH]),.Weight_19(Wgt_9_319[18:19-`WGT_WIDTH]),.Weight_20(Wgt_9_335[18:19-`WGT_WIDTH]),.Weight_21(Wgt_9_351[18:19-`WGT_WIDTH]),.Weight_22(Wgt_9_367[18:19-`WGT_WIDTH]),.Weight_23(Wgt_9_383[18:19-`WGT_WIDTH]),.Weight_24(Wgt_9_399[18:19-`WGT_WIDTH]),.Weight_25(Wgt_9_415[18:19-`WGT_WIDTH]),.Weight_26(Wgt_9_431[18:19-`WGT_WIDTH]),.Weight_27(Wgt_9_447[18:19-`WGT_WIDTH]),.Weight_28(Wgt_9_463[18:19-`WGT_WIDTH]),.Weight_29(Wgt_9_479[18:19-`WGT_WIDTH]),.Weight_30(Wgt_9_495[18:19-`WGT_WIDTH]),.Weight_31(Wgt_9_511[18:19-`WGT_WIDTH]),.Weight_32(Wgt_9_527[18:19-`WGT_WIDTH]),.Weight_33(Wgt_9_543[18:19-`WGT_WIDTH]),.Weight_34(Wgt_9_559[18:19-`WGT_WIDTH]),.Weight_35(Wgt_9_575[18:19-`WGT_WIDTH]),.Weight_36(Wgt_9_591[18:19-`WGT_WIDTH]),.Weight_37(Wgt_9_607[18:19-`WGT_WIDTH]),.Weight_38(Wgt_9_623[18:19-`WGT_WIDTH]),.Weight_39(Wgt_9_639[18:19-`WGT_WIDTH]),.Weight_40(Wgt_9_655[18:19-`WGT_WIDTH]),.Weight_41(Wgt_9_671[18:19-`WGT_WIDTH]),.Weight_42(Wgt_9_687[18:19-`WGT_WIDTH]),.Weight_43(Wgt_9_703[18:19-`WGT_WIDTH]),.Weight_44(Wgt_9_719[18:19-`WGT_WIDTH]),.Weight_45(Wgt_9_735[18:19-`WGT_WIDTH]),.Weight_46(Wgt_9_751[18:19-`WGT_WIDTH]),.Weight_47(Wgt_9_767[18:19-`WGT_WIDTH]),.Weight_48(Wgt_9_783[18:19-`WGT_WIDTH]),.Weight_49(`WGT_WIDTH'b0),.Weight_Select(select_count),.Selected_Weight(weight9_15));
wire [25:0] out_n9;
Neuron neuron_9(.Weight_0(weight9_0),.Weight_1(weight9_1),.Weight_2(weight9_2),.Weight_3(weight9_3),.Weight_4(weight9_4),.Weight_5(weight9_5),.Weight_6(weight9_6),.Weight_7(weight9_7),.Weight_8(weight9_8),.Weight_9(weight9_9),.Weight_10(weight9_10),.Weight_11(weight9_11),.Weight_12(weight9_12),.Weight_13(weight9_13),.Weight_14(weight9_14),.Weight_15(weight9_15),.Pixel_0(pixel9_0),.Pixel_1(pixel9_1),.Pixel_2(pixel9_2),.Pixel_3(pixel9_3),.Pixel_4(pixel9_4),.Pixel_5(pixel9_5),.Pixel_6(pixel9_6),.Pixel_7(pixel9_7),.Pixel_8(pixel9_8),.Pixel_9(pixel9_9),.Pixel_10(pixel9_10),.Pixel_11(pixel9_11),.Pixel_12(pixel9_12),.Pixel_13(pixel9_13),.Pixel_14(pixel9_14),.Pixel_15(pixel9_15),.Clk(clk),.Neuron_Reset(neuron_reset_r),.Out(out_n9));

reg ready_r; // ready register for computation after input is valid
// clock triggered logic
always @ (posedge clk) begin
    // reset at GlobalResetn
    if (GlobalResetn) begin
        neuron_en_r <= 0; // neuron enable set to 0
        neuron_reset_r <= 1; // reset neuron 
        max_en_r <= 0; // disable max select
		max_reset_r <= 1; // reset max select
        ready_r <= 0;
    end
    // reset when Input_Valid goes high 
    else if (Input_Valid && ~neuron_en_r) begin
        if (~ready_r) begin
            neuron_en_r <= 0; // neuron enable set to 0
            neuron_reset_r <= 1; // reset neuron 
            max_en_r <= 0; // disable max select
            max_reset_r <= 1; // reset max select
            select_count <= 0; // counter set to 0    
            ready_r <= 1;
        end
        // wait 1 cycle after input_valid then enable neuron
        else if (ready_r) begin
            neuron_reset_r <= 0; // disable reset
            neuron_en_r <= 1; // enabling the neuron
            ready_r <= 0;  
        end
    end
    // now computation begins
    else if (neuron_en_r) begin
        if (select_count < 60) begin // begin feeding all inputs to neuron
            select_count <= select_count + 1;
        end
        else begin // done with computation, now select max
            neuron_en_r <= 0; 
			max_reset_r <= 0;
            max_en_r <= 1;
        end
    end
end
    //
    // if (Input_Valid || GlobalResetn) begin
    //     neuron_en_r <= 0; // neuron enable set to 0
    //     neuron_reset_r <= 1; // reset neuron 
    //     max_en_r <= 0; // disable max select
	// 	max_reset_r <= 1; // reset max select
    // end 
    // // enable neuron at negedge of Input_Valid
    // if (~Input_Valid && ~neuron_en_r) begin
    //     neuron_reset_r <= 0; // disable reset
    //     neuron_en_r <= 1; // enabling the neuron
    //     select_count <= 0; // counter set to 0
    // end
    // // computation enabled
    // else if (neuron_en_r) begin
    //     if (select_count < 60) begin // begin feeding all inputs to neuron
    //         select_count <= select_count + 1;
    //     end
    //     else begin // done with computation, now select max
    //         neuron_en_r <= 0; 
	// 		max_reset_r <= 0;
    //         max_en_r <= 1;
    //     end
    // end
    //


// max selector
MaxSelect maxselect(
    .clk(clk),
    .in0(out_n0),
    .in1(out_n1),
    .in2(out_n2),
    .in3(out_n3),
    .in4(out_n4),
    .in5(out_n5),
    .in6(out_n6),
    .in7(out_n7),
    .in8(out_n8),
    .in9(out_n9),
    .max_en(max_en_r),
	.max_reset(max_reset_r),
    .max(Image_Number),
    .max_ready(Output_Valid)
);

endmodule
